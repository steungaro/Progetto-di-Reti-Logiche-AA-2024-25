-- TB EXAMPLE PFRL 2024-2025 -- RUAN HUIJUN
 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
 
entity tb2425 is
end tb2425;
 
architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
 
    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");
 
    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 32759;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      1,                                                        -- S
                                                      0, -1, 8, 0, -8, 1, 0, 1, -9, 45, 3, -45, 9, -1           -- C1-C14
                                                      );
    signal scenario_input : scenario_type := (93, 52, 76, -35, 17, 69, -83, -61, 52, 123, -126, 114, 2, 78, -78, 51, -80, 22, -124, -90, 112, 48, -66, 126, -16, -121, -91, 11, -79, 103, 45, -114, 27, -6, -21, -83, -65, 24, -16, 115, 20, -14, 101, -106, -64, -105, 73, -16, 46, 77, 22, 30, -3, 85, 29, 110, 92, 66, -7, -115, 42, -90, -101, -59, 32, 7, -14, 96, -97, 99, 83, 51, -43, 57, 74, 22, 80, 19, -122, -2, -31, 29, -99, 94, -14, 58, 76, -50, -4, -59, -36, -90, -20, -9, -20, -116, 126, 94, 108, -98, 65, 64, 81, -105, -7, 27, 45, -55, -81, 51, 72, 16, -48, 101, -18, 66, 31, -69, -111, -101, 0, -19, -62, 108, 100, 46, 121, 99, 12, 101, -127, -50, 37, 82, -27, -98, -18, -110, -24, 29, 69, -80, -83, -106, -107, 27, 88, 52, 86, 105, 79, -41, -42, -111, -61, -69, 63, -68, -98, -52, -94, -97, 26, 71, 113, 127, 102, -33, -111, -50, 124, 86, -2, -87, 108, 19, 69, 69, -57, 27, 46, -106, 114, -123, -88, -74, -64, 103, -14, -34, -77, 20, -3, 77, -36, -18, 76, -62, 78, 93, 16, 74, 52, -114, 116, 32, 33, 57, -27, 104, -44, -108, 126, -57, -103, -90, -3, -39, -114, 111, 55, -63, 4, -76, -113, 96, 34, 91, -94, -16, 57, 50, -69, -19, 64, -81, -115, -31, 104, -13, -55, -68, 7, -57, 3, 32, -18, -128, 121, -4, 112, 48, 61, -12, 100, 76, -44, 6, 40, -10, 119, -31, -88, -78, 78, 104, -31, 91, -55, -55, -50, 18, 5, 85, 89, -119, -11, -57, -119, -18, 67, 121, -98, 1, -19, -126, -51, 65, 9, 117, -73, 0, -42, -33, 50, -92, -57, -109, -128, 16, -36, -50, -94, 97, -92, 124, 106, 25, -61, 116, -120, -121, 109, -90, 8, -37, -87, 85, -100, 50, 75, -44, -78, -95, 51, 100, -58, 123, 119, -58, 11, -45, 20, 46, -76, 56, 42, -97, -46, 109, -109, -38, 116, -128, 0, -4, -37, 41, -46, -8, -37, -99, 76, 13, -66, -1, -15, 4, -6, -24, 74, -122, 59, -33, 52, 112, -105, -34, -113, -23, -53, -94, 67, -64, -94, -60, 60, -2, 109, -114, 118, -55, -85, 66, 86, -22, -63, -56, 110, 60, 48, 57, 66, -20, -104, -10, -36, -81, 84, -21, 25, -97, 13, -36, -33, 47, 32, -100, -83, 14, -86, -93, 87, -42, 101, 45, 64, -89, 117, 46, 99, 38, -25, 37, -110, -1, -101, -18, 47, 111, 89, -56, -114, -26, 36, -18, -107, -59, 10, -61, 83, 52, -26, 42, -118, -52, -41, 74, -13, -51, -7, -42, 115, 96, 123, -123, -32, -106, -13, -113, -123, -52, -41, -109, 50, 123, 1, 71, -64, -117, -118, -109, 64, -15, 61, 74, 61, -107, 21, -80, -30, -114, 6, -43, 110, 1, -38, -50, 23, 77, -35, 28, -103, 52, 47, 75, 48, -79, 18, 112, -68, 29, -124, 124, -114, 65, 71, 75, 86, -36, 123, -72, -22, 1, 13, -40, -126, 103, 39, 25, 52, -124, -75, 77, 57, 100, 24, -23, -107, -85, -39, -46, 72, -35, -50, 86, -97, -107, 33, 117, -15, 28, -82, 91, -99, 59, -76, -97, 35, 91, 56, -41, 95, 109, -91, 24, 81, 61, -127, 103, 104, -37, -71, 48, 56, 7, 6, 87, 29, -89, 77, -114, 67, 123, 106, 96, 54, -98, 127, -39, 121, 55, 49, 88, 36, 86, -15, -10, 19, -14, -35, -4, 77, 22, -84, 6, -99, 51, -35, 58, 90, -86, 73, 30, -91, 51, -2, 92, 81, -2, -75, 74, -75, 102, 34, 90, 60, -109, -48, -48, 6, 45, 76, -45, -61, 120, 89, -32, 43, -73, -101, 6, -31, 100, -92, 7, 23, 34, -29, -24, -96, 24, -78, -42, -1, 84, -80, -69, 104, 0, 11, -18, -83, -41, 65, -16, -48, 27, 80, 123, 82, 107, 1, -77, 79, 37, 58, -26, -56, -99, 78, -24, 54, -128, 62, -75, 85, 110, -16, 61, -18, 124, -85, 27, -45, 108, -117, 35, 7, 92, 31, -39, 71, -96, 13, 23, 70, -57, 125, -114, -27, 76, -10, -101, 76, -75, -48, 33, -93, 64, -34, 18, 60, 9, -83, -112, -10, -71, 51, 125, -107, -46, -41, 92, -13, 100, -13, -71, -85, -15, -57, 16, -67, 61, 43, -119, 114, 123, 43, -106, 60, -119, 40, -8, 19, 85, 8, -119, -114, -68, -122, -93, 14, -35, -128, -127, -63, -13, -70, -19, 100, 1, 125, -95, -65, 41, -85, -79, 36, 86, -57, -32, 95, 111, 89, -14, 69, -31, -5, 83, 29, 2, 119, -84, 95, 119, -83, -95, -22, -24, 14, -49, 105, 11, -16, -88, -76, 27, -38, 89, -15, 33, -71, -47, 17, -110, 67, -42, -12, -65, -87, -111, 65, -96, -67, 32, -105, -21, 65, 2, 83, -49, 81, 60, 91, -63, 101, -113, 93, -65, 104, -50, 96, -94, 31, -15, -76, -29, 71, 40, 34, 113, 58, -29, -111, 119, -125, -87, -30, 69, 43, -75, -108, -4, 114, 111, 61, 87, 127, 26, -106, 103, 105, 118, -119, 8, -24, -66, 107, -81, 102, 13, -96, 32, 112, -78, 24, 116, -37, 122, 57, -122, -80, 77, 2, -94, 61, -65, 121, 60, 90, -113, 35, 67, -123, 45, -53, -19, 107, -73, 29, 81, 68, 61, -14, 53, 111, -118, 41, -54, -124, -30, -48, -76, -81, 82, -42, 108, -110, -49, 40, 108, -34, -52, 47, -28, 121, 122, 81, 100, -79, -18, 53, 118, -84, -89, 43, -101, -79, -44, -26, -74, 54, 54, -22, 101, 9, 65, 82, 27, -112, -6, 7, -17, 70, -74, 83, 63, -80, 36, 35, -30, -109, -39, -40, -65, 0, -125, -38, 50, -41, 64, 104, -115, -9, -46, 114, -128, -109, 68, 27, -92, -65, -94, 19, -123, -40, -26, 69, 8, -118, -24, 106, -99, 65, -62, -36, -62, -59, 55, 116, 28, -9, 92, 41, 110, -82, 28, 110, -62, -32, 9, -26, 31, 43, 121, 37, -125, -33, -22, 12, -23, 82, -10, 7, 20, 57, 99, 86, 126, 26, 74, 27, -110, 38, -60, -128, 84, 96, 111, -106, -63, -8, -4, 96, -92, -11, 5, -89, 84, 111, 51, -66, 66, -86, 69, -42, 99, 40, -84, 97, -61, 118, -4, -43, 28, 65, -43, -16, 33, -60, 7, 98, 61, -125, 67, 97, -7, -56, -120, -51, -72, 60, 11, 122, 102, -48, -48, 73, 121, -4, 42, -68, -14, -89, 17, -114, 104, 102, -2, 9, -85, -123, -20, 104, -119, -81, 73, 2, -9, 81, 79, 47, 13, -37, 41, -13, 43, 121, -68, 36, -11, 103, 96, 103, -114, -15, 117, 118, -40, -12, -1, 3, -7, 107, -21, 2, -102, -76, -124, 18, -123, 84, -63, 19, -81, 107, -122, 90, 100, -61, -1, -38, -86, -33, -63, -72, 81, -73, -82, -87, 43, 45, 44, -92, 25, -105, 39, 51, -53, 43, -59, -48, -1, 7, 99, 46, -14, 106, 9, -42, -83, -120, 48, -41, -25, 114, 15, -72, -87, 61, -31, 84, -22, -115, 120, -125, -92, 31, 55, -17, -53, 124, 64, 74, 3, 35, -7, 117, 13, -126, -52, 58, -118, 124, -111, -15, 110, 32, 42, -105, -35, -117, 107, 72, -103, 100, 75, -67, 3, 2, 45, 78, -1, -19, 25, -126, -112, -110, 120, 30, -108, -60, -40, -98, -64, -22, 15, -81, -118, -71, -58, -24, -59, -78, -80, -34, -106, 123, 27, 25, -2, -56, -24, 125, 53, -127, 127, 70, -109, 119, -28, -89, -69, 60, -59, -4, -90, 84, 43, -79, -114, 113, 25, -45, -93, 73, 49, -71, 68, -52, 83, -62, 21, -69, -65, -54, -68, -65, -112, -49, -74, -12, -10, -14, -79, 59, 110, -41, 15, 25, 8, 29, 10, -95, 112, 46, 106, 33, 103, 47, 110, 58, 113, 3, 117, -79, 77, -79, -16, 94, 0, 38, -46, 118, -104, 3, 49, -122, 91, -63, 31, -29, 94, -86, 5, 79, 88, -17, -16, 63, -98, -34, -6, -112, 97, -17, -63, 47, 33, 49, 13, -95, -41, 95, -104, -16, -29, 73, -10, -66, -118, -106, 33, 105, -64, -90, 56, -104, 22, -88, 87, 52, 7, -47, 68, -24, 65, -123, -105, -30, 54, 36, 3, -114, 4, 27, -2, 103, -27, 116, -91, -17, -118, 70, -40, -54, 109, -112, -30, 3, -71, -70, -73, 64, 11, 124, -88, -52, -127, -64, 46, 56, 100, -78, 70, -24, 77, -60, -49, -78, -72, -12, 34, -61, -69, 122, 13, -88, -117, 112, 43, -60, -86, 98, -124, 53, 94, -84, -126, 96, -20, 48, 24, -47, 98, -34, 57, 48, 34, -119, 98, 90, -3, 4, -99, 56, -1, 43, 96, 10, 27, 11, 78, 69, -18, 82, -6, -52, 126, -4, -84, -21, -83, 68, 60, -113, -94, -11, 63, 68, -2, 34, 31, 124, -90, 60, 52, 37, -25, 21, -81, -126, -96, 125, 71, 14, 79, -62, 91, 78, 62, -121, -71, 107, 76, 117, 123, 110, -22, 58, 51, 105, -36, -46, 101, 3, -114, 25, -88, -10, -82, -40, -8, -49, -43, -64, 93, -91, 2, 56, 115, -64, 64, -84, -84, 12, -95, -89, -6, 11, 97, -83, -12, -66, -1, -39, 65, 14, 115, 105, -124, -95, -63, -4, -16, 23, 60, -50, 60, -66, -122, 47, -1, 70, 91, 43, -46, 124, 82, 77, 7, 51, 122, 124, 113, -6, -43, 50, -120, -56, 28, -116, -22, 93, 8, 90, -12, -59, -88, -80, 3, -81, 95, -126, 117, 58, 45, -56, 54, -1, -107, -66, -77, -113, -70, -92, 9, 15, 87, 17, 88, -13, 29, -62, -48, -90, -100, 69, -21, -59, 117, 110, -12, 85, 113, -23, 15, 30, 49, -58, -98, 70, 4, -47, 86, 62, -11, -33, -51, -52, 113, -91, 63, 14, -25, -112, 52, 4, 85, -97, 73, 74, -114, -67, 31, 127, 38, -81, 29, -40, -11, 59, -98, 121, -116, 116, 55, 2, -44, -124, 78, -59, -86, 14, 83, 17, 30, 8, -107, -13, 39, 94, -67, 53, -101, 93, 52, 66, -116, -46, -102, 1, -115, -72, -6, -102, -83, -79, 28, 1, -75, -22, 70, -33, 120, 25, 113, 22, -95, -122, -119, 73, 101, -57, -2, -128, -92, -77, 66, -80, 5, 92, 49, 18, -107, -85, 44, -62, -36, -56, 67, 17, 51, 9, 113, 43, -94, 98, -62, -60, 104, -53, -115, 77, 18, 11, 78, 54, 62, 16, 102, -61, -19, 23, 86, 2, 66, 2, 68, -98, 75, 7, 48, -2, -112, 33, -87, -78, 3, -21, -10, -21, 55, 3, -71, -55, -113, -121, -128, 77, 23, 102, -111, -124, -2, 103, 6, -64, -23, -54, -33, -76, 81, -113, 50, 97, 48, 92, -108, -77, -57, 10, 30, 126, -114, 87, -56, -99, 94, -56, 106, -10, -82, 123, -6, 44, 98, -127, 109, -52, -53, -52, 0, -99, -37, -77, 126, -117, -113, -110, -66, -42, 29, 92, -43, 43, 52, 29, 72, 18, 101, 50, -120, -109, 46, 3, 64, 16, 4, 45, 92, 79, 121, -35, 108, -44, 16, 107, -33, 31, 125, 29, 117, 26, -7, -54, -59, -83, 103, -115, 64, 76, 64, 72, 96, -18, -53, 32, 126, 79, -51, 91, 31, -58, -72, 11, 26, 72, -10, 121, -25, -12, 22, -36, -114, -113, 39, -44, -67, 14, -31, 125, -37, -95, 69, -69, 15, -111, 91, 14, 96, -88, -23, -1, -18, 33, -117, -120, -23, 1, -127, 80, 117, 23, -84, -124, 38, 83, -40, 99, -30, 57, 96, 61, 91, 38, 120, -22, 55, 83, 120, 23, 123, -31, -105, -23, -126, -94, -15, -21, 35, -14, -69, 25, -119, -24, 29, 47, -69, 117, 19, 29, 46, -13, -38, 9, -103, -46, 116, 80, -91, 108, -24, -96, -50, -1, 9, -48, 33, 122, 60, -60, -20, 119, 93, -11, -33, -6, -91, 27, -17, 56, -72, -98, -85, 19, 39, -59, 101, 27, -107, -117, 8, -3, -85, 86, 124, 53, -90, 29, 47, 98, 98, -100, 90, 63, 17, -71, -70, 54, 84, 41, -18, -115, 71, 26, 32, -17, 95, 5, -118, 116, 16, 18, -14, 60, -24, -18, -15, 15, -116, -96, -15, 110, -68, -53, 45, 78, 5, 103, 4, -39, 17, 115, -26, -40, 13, -122, 71, -20, 12, 82, -32, -100, -28, 82, 88, 77, -63, -55, -36, -51, -22, 77, -69, 38, -103, 104, -12, 30, 80, 121, 119, -31, 108, -34, 57, -7, -28, 1, 101, 112, -45, -59, -115, 55, -104, 101, 4, -39, -81, 96, 38, 25, 46, 97, -65, 71, 73, 52, -27, 25, 45, -36, 122, 25, 58, 52, -110, -97, -75, 119, -113, 8, -68, -100, -65, -44, -126, 68, 45, -79, 36, -45, 74, -46, -76, -119, -103, 126, 61, -2, 23, -22, 91, 18, -125, 21, -58, -107, 52, -5, -116, 68, -125, -55, 96, -62, 29, 98, -122, -53, -109, 43, 30, 93, 125, 83, 103, -105, 81, 36, 21, -24, -113, -16, 122, -110, -122, -64, -88, 58, 59, -76, -2, 62, -3, -33, -127, -101, -63, -121, -26, -43, 50, -124, -78, 48, 87, -103, 71, 40, 62, -36, -111, 77, 77, -117, 95, 83, -52, -121, 13, -121, -68, -116, 70, 57, -21, 71, 84, 44, 78, -70, -127, 1, -65, -76, -79, -106, -51, 120, 63, -117, -44, 80, 88, -95, 91, 56, 116, -89, 63, 2, -81, 123, 14, 117, 53, 121, 60, 9, 37, 10, 68, 39, -117, -125, 91, -68, -103, -88, -76, 88, -76, 9, 40, -116, 42, 4, 68, 31, 43, 4, -95, 90, -1, 47, 79, -76, 40, 11, 62, -51, -106, 2, 116, -95, 5, 79, -34, 30, 120, 18, -9, -84, -101, -97, -72, 70, 35, 125, -27, -49, 1, 6, -87, -128, -75, 121, -75, 93, 4, 115, -86, 26, -11, -97, 60, 122, 110, -102, 24, 102, 44, -113, -110, 72, -81, -53, 14, 82, -56, 115, -95, 73, -7, -53, 73, 46, -60, 126, 11, 72, 113, 53, -29, -26, 84, -97, -32, 67, -71, 121, 41, 101, -120, 60, 45, -73, -121, -69, -118, -49, -82, -85, -104, 39, -10, 97, -43, 58, 96, 96, 3, 81, 22, 102, -72, -22, -123, 24, -83, -66, 17, 87, -93, 26, 19, 81, 81, 26, -116, 91, 105, -69, -121, -127, 98, -3, 98, -72, -72, 66, -104, 59, 20, 46, 33, 76, -103, 38, -28, -58, 100, 118, -99, -121, 16, 48, 88, -31, -54, 101, -67, -77, -96, -60, -76, -126, 65, -105, -70, 121, 89, -45, 52, -19, -127, -43, -71, -102, 123, 30, -31, 95, 20, -2, 103, -92, -81, 63, 5, -7, 36, 66, 45, 68, -122, 97, 71, 72, 120, -127, 65, 82, -44, -10, -65, -42, 75, -7, -16, 71, -105, 81, 38, 43, -48, 13, 79, -1, -51, -44, 120, 113, -105, 37, 54, -99, 7, -3, 101, -1, -2, 39, -47, 83, -99, 17, -87, 104, -118, 25, 47, -95, -21, -42, 76, 59, 99, 27, -70, -80, 111, -78, -94, -122, 88, 88, -92, -33, -43, -119, 94, 83, 48, -80, 38, 77, 65, 79, 54, 75, -23, -27, 108, 84, 59, 56, 15, 31, -45, 73, 79, -62, 123, 113, -55, 83, 73, -19, -78, -98, -10, -111, 114, -89, -63, 24, 116, -126, -24, 42, 77, 81, -112, 57, 37, 75, -15, -76, -22, 68, 125, -70, -122, 120, -85, -49, 76, 117, 60, 126, -109, -77, -113, -123, -38, -48, 30, -50, -46, -122, 121, -97, 87, -119, 88, -4, 84, -55, 48, -65, -115, 45, -7, -108, 37, 36, -29, -15, 25, -96, -16, 45, -45, -1, 50, 45, 80, -48, 123, -94, -42, 116, -62, -83, 125, -102, 41, 82, -28, -39, -111, -15, -122, 10, 5, 44, -82, 105, -99, 72, -119, 13, -11, -36, -115, -89, -119, 93, -8, -124, 127, 78, 121, -63, 124, 118, -36, 37, 72, 64, 127, 89, -79, -123, -29, 55, 49, 18, 32, 79, -38, 41, -36, 79, -123, -23, 118, -114, -58, -18, -110, -58, -67, -117, 7, -71, -126, 99, 94, 74, 35, 93, 36, 85, 99, -121, 12, 20, 25, -84, -29, 115, 85, 64, 66, 90, -87, 57, 104, -16, -89, 122, 54, -28, -122, -67, 29, -120, -95, -4, 82, 68, -39, -10, 25, -68, -2, -91, 81, -105, -47, -76, -117, -90, 116, 77, -128, -98, 6, 104, 14, 46, 99, -60, -110, 105, 1, 48, 113, 34, -84, 67, -25, 5, -70, -128, 66, 56, -90, 19, 79, -9, 71, 90, 30, 60, 40, 30, 90, -82, 7, -24, 92, -22, 44, 111, -45, -83, 31, -60, 80, 75, -121, -73, -48, -63, -73, -110, 121, -35, 37, 73, 85, -19, 35, -13, -87, -53, -111, -125, -6, 24, -21, -42, -126, -105, -59, -43, -60, 100, 25, -108, 47, 33, -53, -128, 98, 3, -110, 92, 96, 56, 37, 53, -91, -56, -88, -50, 20, -70, -47, -114, 82, 60, -28, 85, 83, 42, -86, -105, 14, 68, -84, -66, -27, -9, -66, -57, 122, -48, -93, 91, -120, 72, 16, -83, -111, 57, -5, 37, 115, 76, 51, 69, 8, -105, 26, -37, 65, 69, -13, -48, 9, 31, 14, 110, -106, 76, -75, -111, -100, -39, 108, -91, -95, -4, -46, -78, -75, 78, 87, -88, 26, 10, 110, -93, 34, 8, -2, -29, -51, 113, 51, 86, 16, -63, 68, 39, -115, 122, 56, -86, -45, 36, -49, -12, -96, 33, 39, -42, -17, -2, -2, -118, -119, -20, -83, 43, 117, 43, -114, -62, 29, 66, -103, -83, -125, 93, 84, -111, 87, 12, -69, -86, -80, 10, 31, -47, -85, -58, 39, 27, 68, -91, 37, 77, 18, 82, -8, 7, -3, 7, 73, -102, -55, 98, -56, -52, 64, -100, -35, 23, 41, 24, 66, 89, -94, -31, -86, -50, 39, 81, 105, -21, 119, 14, -71, 9, -32, 49, -112, 93, -72, 89, 120, 1, 60, -64, 78, -4, -36, -85, -109, -123, 68, 85, 95, 102, -74, -119, -76, 93, 91, -99, -55, 82, 43, 2, -37, -117, -77, -21, 105, -20, -60, 97, 109, -128, -95, 59, -4, -3, 103, 16, 3, 43, -27, -30, 17, 28, -21, 70, -7, -58, 99, 66, -104, 15, -60, -13, 26, -8, 94, 3, 100, -93, -28, 81, -93, 5, 13, 32, -125, -12, -80, 6, -97, 21, 104, 48, -79, -45, -10, 43, 26, -38, -19, 50, 105, 50, -90, 3, -86, -124, -121, -114, -89, -21, 95, -53, 113, -20, 107, 116, 96, -101, -6, 127, 48, -30, 48, 98, 53, -90, 13, -49, 0, 122, -126, -23, 44, -88, 109, 86, -84, 116, 100, -44, -33, 68, 31, -48, -80, 10, -60, -111, 37, 62, -112, -43, -96, 64, -73, 86, 103, 68, -91, -25, 63, -89, 81, -21, -49, 62, -62, -4, 50, -90, 80, -111, 106, -17, -30, -101, 121, 38, -84, 30, -27, -68, 115, 5, 125, -85, -37, 100, 111, 1, -53, 46, 40, -100, -102, 120, 90, -36, -12, 12, 2, -60, 30, -19, 51, -128, 8, 44, 38, 52, -54, -117, 112, -67, 17, 109, -24, 108, 81, -40, -19, -99, -122, -106, -71, -96, -114, -108, -4, 2, 32, 127, 70, -66, -20, -7, -66, 116, -91, 101, 40, -17, 112, 24, 44, 1, 6, -107, -18, -41, -19, 91, -12, -13, 113, 46, 20, 127, 66, -112, 1, -30, -113, -57, 33, -5, 64, 95, -17, 101, 68, -105, -44, 53, 48, -127, -74, -74, -106, 36, 13, 3, 0, -126, 118, -15, 48, 10, -15, -14, 27, 114, 84, 42, -70, -11, -90, 122, -43, 21, 96, -103, 45, -76, 78, -35, -75, -123, 19, -53, 41, -96, 78, -87, -94, 69, 27, 82, -49, -116, -60, 106, 126, -103, 21, -72, 14, 59, -77, 99, -48, -109, 125, 125, -57, 75, -38, -3, 80, 109, 72, -6, -114, 23, 35, -80, -36, -66, -125, 43, -54, -57, 22, -55, -32, -85, 1, 111, 102, 52, 82, -74, 71, 79, -76, -113, 27, 14, 12, -21, -4, -44, 101, 10, 107, 9, 58, -57, 71, 61, 115, -110, -123, 9, -37, -27, 52, 92, -44, 26, 17, -89, 80, -40, 118, -124, -25, 17, 19, 115, 125, -113, -56, 98, 25, -77, -21, -45, -5, -77, -111, -18, -59, -106, 119, 32, -5, 43, -4, 80, -59, -115, 119, -107, -26, 109, -102, 77, -1, 45, 65, -4, 60, -119, -34, -43, -68, 74, 40, 55, 125, 57, -91, -62, 79, -100, 98, -53, 71, -34, -101, -116, -20, -110, -94, 82, 127, -68, 31, -2, 105, -32, 122, 37, -23, -39, 122, 38, -93, 34, -35, -96, -36, 3, -30, -85, 31, -60, -10, -25, 34, 17, -13, -114, 35, 21, 96, 35, 81, 0, -95, 58, 96, -100, -33, -54, -11, -39, 112, 24, 124, -51, 56, -40, 80, -102, 3, -16, -34, 122, 87, -128, 11, -54, -113, -81, 96, 111, 82, 49, -17, 115, -20, -48, -113, 75, 26, 4, -91, 10, -100, -95, 87, 84, -7, 40, 110, 124, -104, -52, 118, 111, -51, 2, -71, -36, 49, -103, -53, 3, 75, 59, -10, -73, -117, 6, -126, 37, -118, -89, -81, -89, -56, -122, 123, 65, 46, 106, 62, 70, -74, 52, 53, 3, -74, 111, 95, 103, -120, -85, -22, 83, 102, 97, -118, 113, -25, -115, 22, -15, -76, 69, 24, -3, 75, 20, -66, -6, -2, 124, -64, 52, 49, 118, -72, 103, 101, -105, 79, 109, -62, -71, 65, -88, -102, 75, -103, 1, 88, 47, 115, -115, -12, 11, 10, -64, -97, 72, 58, 29, 69, 122, -46, -10, 112, 10, -35, 85, 33, -84, 67, 100, -26, 4, -116, 0, -49, -90, -126, -88, 85, 117, -75, -54, 0, 63, 10, 32, 7, -60, -67, -52, -66, 15, 66, -81, -103, -96, -124, 59, -52, 71, 31, 50, -53, 43, -77, 27, 81, -75, 67, 39, -86, 120, 113, 42, 55, -5, -54, -66, 63, 8, 11, 125, -105, -51, -84, -79, -19, -79, 108, 58, 120, 11, -20, -60, -74, 31, 95, -120, 84, 34, 47, 126, 26, 32, 41, -47, -101, 115, 15, 90, -5, -102, 87, 19, -24, -124, 68, 85, -75, 48, 15, -83, -69, 124, -15, -15, 27, -48, -7, -16, 114, -88, -18, 12, 72, -105, 93, 99, -117, -19, 61, 6, 7, 21, -103, 111, 25, 93, 69, 78, 13, -44, 123, 72, -48, -19, -70, 108, 61, 51, -36, 48, 92, 74, -68, 36, 98, -102, 8, 109, 7, -59, -13, -114, 90, 13, 126, -13, -22, 67, -63, 120, -105, -67, 64, -24, 42, 122, -44, -25, 46, 48, -105, 10, -6, -44, -82, -36, -18, 54, -55, 117, 124, 61, -125, 86, -54, -127, -54, 52, 68, 11, 44, 92, 72, -19, -60, -14, -25, 24, 90, -107, -56, 113, 31, 66, -59, 78, -97, 51, 4, -24, 40, 0, -91, 44, -41, -17, 45, 33, -92, -14, -84, 80, -50, 117, -67, 18, -25, 37, -86, -63, 58, -14, -77, -38, -76, -8, -88, -45, -84, 44, 60, 84, -83, 97, 0, 4, -47, -82, -91, -11, 32, -47, -59, 110, -58, 3, 0, 46, -88, 42, 111, 98, -100, -94, -68, -48, 27, -28, 36, 71, -111, -32, 27, -66, -63, -100, 66, 18, -54, 103, -121, 106, -72, -51, 88, -1, 80, -40, -83, 120, -126, -100, 90, -98, -65, -105, -18, 90, -5, -110, 33, 12, -14, -68, 74, 52, -40, 12, -58, 34, -13, -50, 12, 44, 27, -28, -85, -21, 60, -40, -29, 62, -12, -67, 92, 51, -44, -53, 13, 80, -35, -82, -36, 80, -21, -89, 4, 67, 51, 74, -26, -89, -104, 114, 83, 51, -41, 126, -98, -109, -42, 1, 82, 74, 63, 46, -2, -109, 121, -117, 99, -41, -70, -64, -89, 37, -25, 43, -24, -102, -11, 78, -63, 14, 65, -108, -63, -104, -110, -32, -85, -24, 97, 125, -77, 32, 44, 49, 52, 37, 60, 23, 124, 118, 87, -93, 27, -66, 78, -124, -39, -60, 82, 26, 82, 19, 47, -109, 43, 65, -13, 87, -86, -43, 84, -35, 117, 0, -114, 41, -90, 74, -63, -94, 65, -104, -58, -36, -41, -108, -32, 48, -40, -77, -54, -86, 70, 121, -66, -14, 59, 49, -55, 101, -122, -99, -62, 124, 30, -48, 37, 68, -102, 102, 102, 91, 127, -84, -72, -42, -63, 24, -122, 25, 75, -48, 68, 18, -54, -126, -124, -123, 51, -51, 106, 58, -22, -84, 54, -120, -4, -37, 76, 22, -62, 51, -14, -63, 95, 42, 23, -96, -62, 29, 58, -114, 109, -2, 32, -73, 0, 36, -68, -77, 113, -90, 109, -37, -46, 35, -28, 78, 127, -80, -27, -63, 99, 87, 2, 67, 1, -103, 99, 67, 54, 29, 81, 35, -101, -15, 91, 27, -107, -105, 79, -122, -66, 60, -30, 16, -32, 70, -33, -33, 118, 68, 32, 90, 27, -94, 29, -100, -69, 0, 95, 113, -98, 49, 20, -71, -94, -17, 85, -72, 7, 36, -66, 69, -32, 32, -43, 64, -26, 52, -97, -35, -8, 63, -73, -109, 97, 84, -81, -100, -44, -113, -115, -14, 64, 34, 44, 98, -111, 1, -102, 24, -91, -39, -35, 5, 121, 51, -58, -32, -25, -27, 61, 96, -91, 116, 115, -122, 72, -93, -93, -100, -78, -80, 15, 114, 82, -69, 84, 100, 60, 111, -4, 97, -56, 90, -26, -63, 13, 44, 33, 116, -110, -34, 84, -73, -46, 72, -67, -102, 107, -32, -73, -99, 17, 70, -113, -29, -127, 99, -57, 61, 82, 68, 30, -102, 30, -124, -36, -85, 49, 125, -97, 67, -36, 116, 122, 46, 60, -73, 73, 39, 24, -128, 68, -87, 70, 83, 12, 71, 54, 84, 4, 9, 24, -94, 35, -74, -90, 127, -31, 87, 125, 0, 26, -39, -12, 20, -121, -80, 76, 80, 87, -28, 80, 27, 13, 22, -18, -103, -35, -91, 109, 97, 46, 5, -125, -47, 59, -86, -47, -100, -127, -50, 29, 28, 39, -111, -80, 46, -62, 124, -1, -103, -32, -49, 53, 109, 102, -93, -121, -61, -56, 116, -91, 118, -6, -88, -56, -75, -46, 25, -46, -44, 103, 111, 112, 14, -128, -96, -68, -62, -99, 59, -36, -3, -117, -111, -21, 113, -76, -14, -76, -3, -26, -39, -13, 96, 2, 59, -106, 84, -44, -24, -88, -69, -41, -104, 73, -41, -71, -122, 26, -42, 65, 118, 83, 76, -121, -66, 61, -69, 48, 114, 56, -105, -53, -84, 119, 77, 103, -115, 34, -68, -11, 74, -9, 76, 99, -63, -92, -100, -57, 62, -14, -120, 52, -59, 85, 59, 4, 18, 118, -76, 4, 47, -53, 80, 91, -61, 29, 66, -48, -65, 126, 70, -118, -10, 18, 109, 55, 54, -119, 126, -12, -5, -122, -88, 64, 91, 99, -60, -18, 90, -7, 114, 9, 68, 66, -28, -121, -32, -90, -40, 31, -91, -98, 41, 27, 48, 22, -46, -25, 31, -48, 91, -102, -42, -124, 91, -78, 103, -97, 32, 65, 24, 18, -54, -35, -43, 46, -28, 53, 85, 60, -44, 122, 90, 126, 21, 11, 20, 103, 114, -76, -73, 77, -50, 13, 81, -87, 63, 57, -55, -33, -6, 97, 114, 69, -66, -57, -13, 35, 124, -56, -33, -48, -62, -70, -50, 87, 69, 99, 62, 55, -105, 117, 4, -27, 3, -42, 15, -62, -113, 88, 34, 9, 57, 20, -50, 120, 91, 66, 27, 87, -118, 122, -89, -51, -76, -10, -92, 121, -39, 99, 48, -16, 88, -75, 85, -37, 11, -28, 30, 26, -68, -64, -93, 118, 84, -14, 110, 47, -76, 9, 6, -66, 3, 45, 11, 56, -93, 48, 49, -4, 19, -30, 108, -21, 23, 66, 71, -94, -90, -27, 60, -29, 37, 95, -39, -7, -47, -57, -88, 5, 80, 46, 68, -45, -37, -49, -117, -1, 127, 61, 123, 18, -97, 104, 126, 54, 42, 69, 88, 80, -86, 20, -77, 79, -13, 12, -56, 69, 83, -16, -54, 35, -98, -114, 119, -7, -34, -126, 120, -35, 63, 116, 112, 94, 92, 110, 20, 6, 51, -20, -42, 93, -128, 10, 44, -12, -106, 116, -71, 106, -28, 3, 13, 2, 18, 4, 123, 112, 7, 116, -51, -58, 104, -67, -91, 68, -85, 57, -54, 94, -90, 32, 59, -90, -86, -25, 26, -63, -37, 83, -85, 63, -41, 56, -63, 105, -67, -67, 89, 68, -79, -90, -118, -103, -28, -81, 93, 15, 105, -89, -18, -113, 71, -87, -75, 114, 17, 80, -77, 108, 35, -34, 44, 122, -106, 109, 99, -45, -86, 60, -105, -37, 99, -94, -12, -57, -47, -47, 86, -70, -8, -60, -55, -64, -18, -1, -78, 127, -49, -27, 107, 114, 67, 23, 109, 89, 5, 80, -83, 47, 13, -60, -117, -16, -26, -1, 55, 56, 81, 13, 114, -55, 82, -68, 9, -64, 59, 59, -65, -118, -96, -86, 124, 99, 66, 105, 61, -57, 58, 106, 118, -57, -82, -127, 55, 21, 1, -18, -51, -46, 123, -65, 27, 77, -5, -91, -115, -74, 96, -52, -64, -127, -9, -67, 100, -71, -90, 33, 0, 96, 11, -10, -89, 58, -8, 94, -49, 121, -52, 28, -53, -56, 91, 102, -107, -41, -117, -93, 13, 108, -17, 78, 109, 102, -117, 81, -97, -79, -13, 31, -110, 126, -106, -71, 56, 14, -104, -121, 7, -28, 35, 82, 44, -1, 56, 66, 86, 68, 101, -29, 48, -44, -79, 29, -69, -68, -18, -38, -18, 97, 122, 0, 96, -112, 57, 24, 30, 81, 32, -91, -74, -61, 119, 98, 66, 47, 36, 24, -13, 9, 124, -93, 94, -83, 64, -103, -22, -81, -13, 88, -112, -19, -40, 112, -3, -111, 9, -101, 99, -87, -64, -103, -20, -73, 123, -81, 103, 32, 71, -38, -87, 67, -2, -121, 113, -66, -96, -37, -19, 20, -77, -2, -127, 11, -18, -1, 28, 119, 26, -1, -96, 91, 24, 13, -110, 20, 60, 121, -76, 3, -44, -35, -57, 82, -27, -72, -112, 5, 19, -2, -103, 70, 124, -101, -47, -22, 26, 109, -30, -76, -19, 2, -113, -123, -113, -94, 25, 75, -101, 77, -49, -17, -85, 22, -63, 16, 78, -46, -107, -31, 80, -81, -89, 76, -54, -8, -74, 100, -27, 24, -104, 82, -101, -88, 88, -86, -54, -15, 118, -27, -65, -59, 85, -22, 91, -106, 122, 41, -24, -113, -118, -72, -66, -79, -124, 8, 41, -69, -20, -114, 83, 5, 97, 110, 45, 57, -103, 119, -86, -113, -36, -23, -44, -79, 83, -81, -56, 77, 88, 48, 93, 98, 105, -101, -109, 109, 36, 60, -88, -112, 74, 124, 21, 43, 106, -62, -28, -125, -71, 15, -110, 22, 120, -26, 71, 76, 21, -113, 25, -19, 64, -10, -49, 41, 18, -30, 22, -74, -98, 63, -58, 105, 59, 92, 20, 37, -98, 121, 41, -40, 8, 59, 110, 0, -94, 53, -52, 55, 69, 102, -91, 5, -36, -12, -82, 110, 87, 68, -92, 117, 3, -21, 94, -66, -57, -13, 100, -27, -20, 13, 61, 116, -56, 43, -12, -22, -31, 65, -94, -90, 39, -57, 43, -125, 59, 89, 114, 18, 29, -106, 8, -95, 1, -26, -33, 72, 89, -61, -82, -59, 80, 107, -71, -103, 23, 46, 3, 120, -17, 37, -98, -106, 108, 73, -103, 40, 34, -117, -70, -65, -94, 66, -32, 35, -87, 64, -20, -126, -125, 26, -56, 84, 5, 1, 109, -100, -81, -16, -108, 30, -106, -78, 52, -126, 123, 78, 42, 29, 89, 101, 93, 123, 39, -67, 31, 80, 125, -117, 83, -127, 37, -101, 85, -86, 28, 66, -57, 76, -78, -37, -22, -56, 14, -97, -53, 9, 109, 117, -89, 70, 90, -124, 66, 2, -63, -31, -46, -65, -20, -91, -64, -111, -64, -107, -69, 93, 87, 2, 41, -119, 94, -109, -46, -20, -78, 29, 117, -97, 18, -100, 102, -19, -96, 40, 111, -30, -119, -63, 33, -11, -25, 97, 6, 39, 118, 65, 4, 77, -60, -83, 86, -94, -63, -88, 14, -13, 69, 3, 19, -40, 32, -7, 69, 64, -95, 52, -94, -86, 117, 67, 31, -36, 36, -91, -124, 26, 102, 8, -25, -86, 54, -66, -52, 119, -26, 90, -22, -84, -34, 125, 4, 126, -10, -55, 62, 23, 125, 97, 65, 114, 36, -32, -49, -55, 5, -45, 99, -20, 91, -53, 22, 17, 9, 99, 8, 111, 61, 115, -101, -101, 112, 31, -103, -25, 104, 88, 126, 101, 57, 64, 88, -35, -96, -89, 38, 38, -6, 10, -110, -43, 85, 40, 103, -34, 11, -17, -51, -55, -30, -23, -28, -45, -120, -2, 58, 113, -42, 56, 86, -113, -8, 46, -20, 25, 85, -109, -65, -49, 29, -47, 37, -14, 121, 12, 80, 5, 123, -99, 78, -34, 6, -78, 49, 15, 48, -21, 0, -122, -93, -42, -107, 28, -123, 2, -75, 90, 21, -12, -86, -78, 69, 79, 36, 62, -37, -12, -61, -42, 17, -111, 52, -104, -60, -27, 39, 116, 80, -89, 123, 116, -3, -112, 16, 2, 18, 69, -35, -89, -71, 7, -39, 126, -42, 125, 60, 49, -15, -128, -121, -125, -111, 60, -101, -43, -95, 66, -54, 114, 105, -59, 102, -26, -43, -10, 105, 104, -69, -58, -113, -12, 77, -23, -14, -93, -26, -82, 84, 88, -82, 91, 91, -64, 23, 118, 21, 57, 56, 95, 43, 33, -92, 17, -121, -6, -121, 112, -30, -62, -74, -15, 54, -125, 90, -88, -90, -63, -42, 122, -103, 5, 86, 116, 69, -19, 106, -38, -90, 34, -70, 81, -61, -34, -30, -54, 88, -23, -69, -70, 43, -15, 44, -31, -11, 6, 9, 27, 71, 96, 22, 96, -27, -20, 84, -86, 89, 62, 4, -128, -32, 62, 81, 35, -99, -76, 110, 117, 29, -87, -80, -55, 26, 92, 42, -113, -30, -76, 43, -86, -108, -63, -118, -7, 45, 95, 35, 6, 29, -89, 6, 126, 102, -40, 33, -125, 12, 15, 120, -87, 56, -88, -14, -45, -124, -99, -30, -25, -47, -115, 17, -27, -50, 27, 94, 123, -6, 1, 2, -104, 40, -120, -106, 14, -32, 55, 17, 108, -57, 10, -106, 127, 50, 8, -46, 55, 37, 53, -98, 118, 66, 47, -37, -111, -54, -71, -116, 69, 58, 14, 93, -29, 23, 115, 113, 119, 42, 3, 100, 113, -115, 122, 113, 63, 2, -61, -10, -88, 120, 20, -98, 59, -61, -6, 76, 14, 51, 88, -45, -18, -25, -80, 81, 126, -93, 66, 117, 77, -59, 89, 63, -46, 83, 48, -110, -42, 115, 8, -2, 108, -99, 28, 39, -32, -106, -13, 110, 74, -53, -63, -72, 50, -15, -119, 48, 20, 75, 38, -30, -111, -1, -95, -29, -45, 81, -11, 41, 68, 126, -89, 48, -101, 67, -41, -5, 90, 74, -22, 36, -106, 43, 92, 72, -99, 101, -7, 49, 48, -97, -109, 65, 30, -76, -91, 113, -123, 26, 26, 74, 24, 65, -6, 51, 5, 82, -81, -33, 28, 25, -125, 50, -60, 95, -5, -31, 68, 116, -109, -12, -109, -90, -74, 49, -37, -37, 35, -32, 117, -67, -86, 14, 127, 37, -63, 4, -9, -16, 99, -109, -119, 102, 70, -50, 69, -63, 47, 9, -75, 66, 125, -56, 105, -77, 121, -60, 14, 28, 36, 4, 90, 79, -110, 89, -12, -45, -35, 107, 68, -64, 126, 77, -90, 68, -101, 107, -123, 75, -12, -70, 13, -15, 2, -10, 37, -4, 58, -77, -104, -33, 55, 114, -82, 73, 75, 34, -99, -88, 13, 97, -24, 11, 46, 14, -48, 74, -7, -43, 21, 109, 16, -94, -33, -110, 25, -124, 14, -45, -73, 39, 50, 111, 25, 96, 56, -27, 2, 85, 13, -113, 54, 118, 27, -27, 4, 107, -81, 126, -64, 68, 107, 80, 102, -54, 99, -1, -50, -15, 83, 6, -104, 5, -11, 50, -26, -83, -105, 104, -125, 36, 120, 57, 26, 19, -98, -97, -2, -51, -99, 62, -111, -120, 15, 120, -45, -14, -9, 33, 99, -54, -89, 124, 80, 28, 46, -74, 74, 69, -98, 77, -23, -106, 6, -124, 41, 37, -93, -89, 114, -64, 102, -124, -56, -11, 124, 27, 103, -13, -67, 74, 62, -28, 70, 14, -127, -12, 68, 75, -71, 98, 24, 35, 121, -98, 39, 34, 67, 74, 74, 54, -118, 48, 58, -46, -91, 54, 110, -116, -87, -85, 86, 103, 15, 29, -11, 16, -111, -71, -37, -53, -100, 115, 110, -107, -110, 21, 55, 85, -33, 1, 11, -23, -79, -59, 59, -42, 123, 41, -30, -91, 84, -71, -116, -28, 86, 2, 116, 103, 59, -48, -78, 87, -61, -96, 108, -43, 53, 36, -85, -108, -91, 54, -3, -41, 124, -71, 45, 119, 98, -112, -100, 55, -55, -87, -101, -97, 43, -113, -122, -26, -33, -71, -66, 35, -39, -86, 120, -113, 78, -93, -93, 116, 90, 33, -53, 86, 90, 120, 77, 60, -120, 106, -13, -47, -109, 14, -16, 62, 30, -9, -92, 125, 48, -30, 32, -119, 13, 25, -104, -37, 60, -68, -49, 22, 93, 26, -20, 55, 19, -70, -13, 27, -92, 103, 109, -73, -11, -35, 117, -109, 84, -103, -111, 4, -4, 49, 14, -119, -54, 38, -28, -121, 98, 52, 29, 63, -50, -118, -10, 97, -60, 106, -3, -24, 81, -22, 31, -58, 71, 20, -38, 28, 45, -21, -96, -87, -100, 46, -78, -25, -43, 23, -18, -73, -53, -117, 119, 25, -107, -19, -5, -39, -41, 120, 65, -88, -30, -32, -17, -87, 116, 73, 69, 34, -76, 102, 75, -48, 20, 126, 55, 105, 21, -91, -95, 96, -79, -104, -7, -58, 5, 116, 32, 93, 108, -31, -123, -50, 66, -12, -8, 54, -67, -67, -40, -15, -93, -92, 66, 56, -94, -7, 33, 55, 31, 66, 23, 80, 90, -112, -106, -32, -123, 54, -67, 113, -104, -62, -64, 90, 55, 56, 16, 116, 117, 105, -26, -103, -115, -88, 81, -81, 33, -14, 102, -64, -75, -3, -112, -113, 13, -89, -17, 18, 93, 44, 4, 117, 111, 68, 79, 38, -4, -32, 26, -15, -55, -128, 10, -42, -88, -37, 5, 74, 78, -21, -118, -125, 104, -101, -110, -11, -62, 2, -120, -97, -82, 12, -107, -99, -48, 100, 67, 76, -60, -34, -67, 13, -34, 72, 99, 7, -93, -24, -47, 113, 83, -37, 116, 59, -10, -121, -79, 56, 9, -71, 88, 55, 69, 109, 85, -107, 81, 24, 97, -106, 118, -98, 35, -43, 102, 7, 92, -118, 111, -83, 123, 67, 8, 112, -2, 127, 119, 47, 55, 0, 104, 15, -73, 45, -4, -116, 66, -50, 37, 35, -28, 27, 66, -121, 112, 40, 14, 76, 50, -2, 121, 46, -63, 2, 30, 63, 1, 21, -17, -72, -107, -41, 72, -52, -123, -60, -39, 71, 18, 126, -21, 118, 25, -83, 126, 10, 85, 12, -42, 8, -118, -48, -74, -53, 82, 84, -117, -45, -23, -6, 11, -2, 81, -45, 74, 86, 24, -93, 30, -86, -95, -119, -95, 59, -74, -97, -59, -117, 43, 27, 19, 54, 107, 73, -127, 61, 29, -116, -112, -122, 6, 28, 4, -40, 111, -49, -82, 7, -14, 76, 50, 20, 85, 83, -49, -117, 114, 20, -105, 29, -81, 42, -45, -101, -12, -43, 88, -111, -31, 105, -104, 104, 5, 28, -64, -12, 107, -18, 124, -34, -69, 46, 114, -112, 1, -63, -100, -13, 85, -77, -112, -124, 93, -28, -97, -47, 57, 120, -29, -102, 97, -5, -126, -26, -105, -62, 90, -125, 49, 86, -31, 108, 4, -45, 124, -123, 20, -104, -8, -23, -53, 9, -19, -87, 109, 13, -6, 38, 5, 93, 64, -26, -40, 67, 76, -16, -123, 38, -13, 54, -3, 84, 34, -127, -89, 31, -121, 59, 55, -1, -92, -125, -120, 17, -84, 117, -98, 38, 27, 35, 4, -36, -119, 92, -97, 85, -52, -92, -4, 63, 91, 121, 19, -3, 122, 58, -100, -127, -11, 84, 1, 25, 87, 9, -85, -125, -1, -55, 41, -102, 109, -83, -10, 118, -118, 21, 76, -42, 58, -56, -106, 21, -63, 41, -110, -69, -28, -81, -67, 89, -125, 62, -13, 90, -57, 30, 93, 70, 103, 6, 97, 84, 52, -41, 75, 62, 109, 23, -108, 39, 95, -86, -68, -96, 84, -50, -37, -72, -3, 24, -111, 0, -42, 4, -38, 30, -94, -73, -28, -118, 62, -59, 94, -14, 29, 41, -80, 10, -64, -60, -79, -97, -17, -19, -65, -61, 59, 27, -5, -71, -77, 12, 57, 10, -111, -108, -88, -77, -53, 12, -67, -119, 82, -100, -5, -17, 69, 43, 121, -122, 112, -86, -91, -33, 23, -27, 34, -46, -128, -99, 11, -77, 41, -59, 61, 58, -39, 101, 110, 36, -14, -85, 46, -60, -57, -87, 51, -115, 85, 44, -109, 69, 86, -72, -92, -19, 29, 70, 63, 29, 99, -53, 81, 12, 16, 14, -57, 105, -12, -75, 13, 102, -32, -69, -86, 40, -27, 93, 53, -70, 9, 72, 127, -33, -128, -93, 76, 30, 105, 11, -69, 76, 86, -116, -40, -26, 27, 31, -49, -113, 84, 93, 117, -75, -104, -97, 93, -3, 124, 18, 55, 5, -38, 54, 100, -38, 89, 48, 120, 66, -69, -76, 14, -110, -64, 103, -8, 91, 6, 72, 106, -37, 37, 95, 16, 61, 126, -19, -69, 122, 127, 114, -1, -39, 41, -29, 51, 2, -109, 44, -59, -49, 96, 83, -31, -96, 58, 89, 124, -63, 33, 102, 28, -58, 70, -84, -124, 68, 25, -65, 63, 24, -79, -66, 113, 90, 34, 36, -35, 53, -48, 34, -124, -80, -11, -27, -47, -80, -65, -51, -15, 96, -77, -115, -89, 121, -71, -85, 62, 82, -22, -3, -22, 27, 59, -37, -10, -35, 127, 83, -109, -48, -11, -105, 0, 106, -3, 81, -102, 60, -98, 11, 28, -46, 24, 67, -53, 81, 110, -119, 35, -40, 6, -115, 116, -62, -24, -22, 31, -24, -67, 50, 56, 50, 74, -72, 28, -57, -118, 55, -125, -88, -62, 31, -6, 91, -29, 70, 44, -47, 79, -48, 42, -42, -35, 30, 24, 70, -120, -73, -82, -59, 106, 102, 119, 52, -98, 19, 123, -88, -54, 126, -47, 13, 29, 75, -24, -128, 17, -108, -46, -31, -28, 124, 55, 66, 26, -49, 8, 34, 6, 54, 103, -16, 28, 94, -92, 58, -15, -97, 99, 60, -99, -76, -55, 59, 127, 49, 59, 17, 69, -115, 114, -86, -119, 41, 108, 35, 120, -12, -59, -2, -86, -84, 111, 70, -118, -109, 0, -4, -77, -29, -72, -48, 23, 1, -117, 23, -78, 71, -88, 119, 84, -102, -95, 94, 67, -115, 1, 59, 1, 71, -71, 43, 115, -88, -15, 126, -68, 114, -6, -17, -43, 50, 63, 109, -77, 75, 4, -27, 18, 44, -36, -26, 70, -2, -60, 9, 11, 70, -60, -115, 13, -3, 56, 0, 38, -86, -2, 98, -100, 120, -47, -15, 42, -112, -34, 93, 91, 98, -62, -19, 14, 31, 84, -44, -99, -104, 93, 40, 94, -95, 53, -21, 31, -18, 108, -59, 24, -22, -89, 52, -29, -8, -91, -115, 8, 4, 107, -28, -26, -83, 81, 117, 76, 37, -55, 105, 62, -89, 18, 28, -56, -57, -120, 103, 53, 116, -84, -51, -34, -45, -127, 65, 75, -89, 79, -44, 43, 58, 56, -111, 103, 9, -122, 52, -81, -48, 29, 109, -9, -81, 9, 63, -9, 17, 39, -84, 5, 83, -6, 100, -89, -5, 37, 114, 34, -12, -58, -51, -82, 126, -33, -106, 8, -27, 74, 55, 53, -25, 36, -84, 23, -83, 108, -114, 63, 19, -70, -60, -26, 52, -88, 13, -80, 78, 0, 82, -62, 70, -96, -15, 69, -1, 7, -51, 100, -47, -124, 26, 56, 40, 70, -49, 85, 50, -35, 20, -59, 24, 89, 44, -52, -127, -71, -4, 79, 57, -49, -110, 0, -17, 3, -59, 110, -118, 18, 82, -37, 22, -20, -109, -66, -77, -29, -109, 101, 64, 40, -85, -40, 1, 87, 37, 2, -112, -95, -46, 74, -16, -28, -54, 95, 103, 15, 77, 113, -95, 32, -52, 55, -116, -33, 117, -65, 66, -120, -91, 3, 48, -48, 91, -79, -89, 0, 52, -73, 34, -122, -127, -110, -22, -53, 114, -47, 90, 63, -62, 123, -33, 14, 50, -20, 109, 39, 43, 48, 48, 80, -77, -32, -96, -114, 18, -57, 15, -58, -1, -79, -52, 0, -61, 54, 76, -75, -121, 38, 117, -55, 34, -44, 87, -44, 64, 68, 124, -20, -12, 44, -68, 39, -116, -35, 54, 30, 36, -59, 100, -93, -10, -80, 36, 57, 102, -16, 111, 109, -106, 100, -74, 56, -72, -115, -115, 121, 82, -119, -27, -58, 53, 33, 110, 65, 126, 36, -32, 35, 105, -60, 70, -33, -11, -22, -104, -37, 90, -121, -55, 113, 107, -1, 41, -92, 13, 54, -99, -33, 63, 2, 37, -12, -93, 19, -74, -94, -73, 22, 69, -96, 90, 11, -1, -49, 118, 24, 43, 80, 31, 116, 65, 11, -13, -21, 47, -128, -95, 76, -33, 97, -50, -123, -43, -15, 24, 11, 19, 80, -95, -40, 112, 124, 100, -16, -53, 90, -120, 118, 42, 39, 106, -20, -78, -34, 87, 97, -34, 120, 45, 62, 89, 123, 67, -81, -19, -37, 58, -128, -85, 92, -39, -100, 88, -67, 12, -93, -105, 20, -102, 65, -69, -124, -83, -18, -30, -124, -49, 65, 125, 125, -1, 86, 120, -62, -123, -27, 29, 64, -26, 73, 28, 63, 101, -12, 124, -15, 23, -109, -123, 49, 84, -64, 54, -126, 46, -104, -122, 126, 89, -125, 123, -40, 90, 115, 26, 95, -39, -72, 31, 63, -127, -69, -2, 102, 47, -6, -41, -57, 13, -36, 120, -31, 28, 46, -29, -53, 71, -22, -55, 32, -19, -60, 121, -57, -73, 19, -89, 16, 75, 70, -49, 76, -126, 77, 50, 49, -57, -119, 120, 84, -27, 113, -74, -126, 31, 25, -51, -26, -125, 22, -121, -15, 90, -128, 56, -111, 19, 95, 34, -33, 38, 113, -85, 40, 63, 94, -39, -122, 103, -46, 91, -51, -61, -111, -49, 98, 42, 28, -55, 46, -78, -48, -97, -116, -48, 87, -99, 99, 55, 63, -62, -35, 49, -18, -123, -16, -52, -34, -10, -77, 48, -47, 0, 115, -30, 79, 86, -115, -21, -97, 59, 29, -17, 90, 41, 63, 49, 71, 34, -24, 6, 101, 69, -73, -45, 74, 39, 31, -87, -98, 82, 89, -17, -45, 77, 82, -94, 35, 95, 14, 66, 26, -85, -79, -12, 85, 112, -91, 28, 18, 14, -94, -9, -45, -38, 74, -98, -127, -23, -57, -97, -68, -96, 15, 15, 109, -31, 49, 16, -64, -65, -46, 90, -21, 3, -50, -64, -13, -13, 92, -122, -127, 126, -3, -43, -40, -56, -13, -38, 49, 58, -7, 109, 90, -120, -4, 72, -23, -82, -40, 41, -19, 43, 3, 88, -82, 81, -104, 34, -59, 116, 40, -58, 115, -91, 27, -53, -19, -114, 37, -97, 72, -97, -116, 35, -89, 9, -21, 17, 55, 67, -70, -92, -18, 62, 125, 29, 15, -107, -65, 84, -118, 103, -101, 125, -116, 54, -56, -6, 69, 110, 25, 13, -115, 37, -80, -76, -82, 27, 69, 101, -33, -128, -118, 77, 62, -121, -22, -51, -100, 41, -94, -90, 16, -67, -93, 29, 115, -20, -105, 56, -38, 48, -58, -25, -43, -10, 27, 4, -110, -31, -23, -15, -31, -13, -66, -97, -6, 41, -20, 23, -46, 14, 61, 99, 75, 97, 0, 63, -51, 23, -9, 39, -57, 61, -114, 28, -76, 41, -96, -58, -118, 10, 55, -21, 125, 117, 10, -8, 30, 119, -113, 113, 5, 76, 84, -47, 45, -44, -112, 122, 107, 7, 33, -78, -59, 47, 78, -7, -39, 111, 63, -29, -7, -10, 79, -10, -21, -39, 110, -118, -48, 125, 123, 86, 74, 79, -89, -9, -93, -73, -14, -114, 62, -109, -64, -125, 67, -114, -4, -100, 125, -69, -1, -10, 49, -50, 109, -99, 40, 91, -89, 120, 89, -94, 78, 35, 113, 117, -102, -108, -84, 12, -94, 107, 32, -30, 110, -29, -16, -21, -1, -18, 38, 126, 100, -40, -51, 81, -11, 117, 45, 28, 109, 6, 62, 60, -87, 47, 49, -61, 67, 94, 80, 101, 73, -16, -57, 55, 83, 55, -94, -46, -91, 73, -48, -118, -95, 29, 91, 22, 18, 8, -78, 0, -114, 112, -68, -73, 31, 109, -5, -30, 75, -53, -57, 20, 59, 14, -52, 14, -59, -18, 96, -21, -73, -80, -11, -40, 78, -48, 110, -32, 89, -96, 96, 103, -112, -100, -97, 47, -118, 26, -111, 85, 101, -40, -22, 32, 102, 54, -82, -84, -92, -114, 23, -36, -66, -116, 52, -116, -36, 35, -19, -75, 67, -51, -99, 84, -22, -68, 3, -12, 86, 21, -55, 59, 109, 51, -37, 84, -23, 9, -128, 14, 23, 23, 106, 85, 35, 30, 98, 127, -63, -49, -75, -123, 28, -46, 89, -122, 14, -36, -6, -28, 113, 68, -97, 95, -9, -6, 51, 97, -125, 51, -17, 26, -54, -39, -17, 109, 119, -47, 108, -71, 32, -95, -66, -67, -13, -105, -61, -127, -13, 62, -27, -27, 2, 4, -60, 121, 126, 119, 90, -127, 42, -55, 27, 116, 34, -117, 97, 26, -36, 77, 83, 125, 111, -111, -70, -30, -88, -3, -28, 27, -69, 73, -128, 61, -50, -60, 55, -52, -69, 17, -50, 101, 91, 105, 89, -3, 116, 58, -105, -47, 8, 106, -50, -9, 123, 8, 89, -93, -123, -67, 63, -63, -121, 63, 126, -43, -124, 53, 33, -65, -57, 111, -91, -94, 89, 126, 31, 77, 57, 55, -98, -63, 33, -20, 56, 29, 116, 17, 64, 122, 79, -1, -69, 86, -65, -71, -85, -61, 111, 76, 2, -74, 60, 39, -40, 21, 38, 119, -30, -33, 46, 1, 32, -48, 109, -40, 109, 98, 105, 45, 92, 56, -83, -105, 14, -20, -48, 57, 47, -65, 6, -79, -11, -62, 89, 77, 87, -1, 69, -71, 94, -13, 58, -2, 67, 40, 86, 48, 10, 63, -34, -26, -8, 11, -3, -122, 119, 77, 64, 38, -115, -58, 87, 2, 8, 48, -48, -33, -81, -107, 24, -115, 8, -45, 11, -52, 123, -31, 124, 5, -95, -38, 107, 25, 101, -24, 31, 92, -75, -33, 2, -62, 37, -38, 69, -83, -118, -107, 12, -70, -86, -91, -57, 50, -8, 83, 126, -13, -76, 123, 120, -43, -43, 99, 110, -69, -53, 14, -105, 0, 109, 26, 67, 19, 116, 8, 64, 126, 29, -51, -72, 71, -14, 0, -7, 106, -45, -8, -35, 7, -13, -43, 93, 72, -72, 75, -125, 3, -39, -101, -125, -57, 53, 70, 90, 41, -50, 26, 39, 107, 103, 96, 50, -39, -32, -84, -61, 51, 36, 32, -70, -105, 117, -105, 95, -83, 99, 99, 48, -68, 126, 52, 3, 51, -6, -35, -36, 73, 120, -125, 52, 95, 99, -25, -71, -61, 19, -4, 118, -73, -99, -79, -50, -110, -56, -83, -64, -85, -112, 112, -24, -114, 36, 107, 65, -97, -55, -99, 104, -63, -95, 28, -96, -124, -125, -39, -56, 22, 86, -66, 77, 115, -17, -101, -123, 56, -55, -59, 99, -39, -74, -53, -24, 90, -73, -87, 121, 0, -57, 97, 65, -24, -2, 97, -20, 1, -69, 52, -104, -111, 115, 101, -124, -30, -127, -119, -102, -54, -49, 126, 35, 5, -55, -117, -33, 0, -75, -39, -128, -4, -70, 65, 100, 56, 35, -48, -70, 94, -123, -46, 111, 120, -73, 115, -38, -72, 124, -11, 2, -53, -13, -90, 80, 60, -79, -80, -67, -26, 9, -67, 98, 67, 127, 70, -4, 34, -105, 54, 0, -100, -120, -17, -108, -65, -30, -18, -8, -34, 99, 122, 42, -42, -96, -6, -109, -46, 42, -48, 56, -77, 13, 27, 119, 12, -31, -13, -82, -8, -87, 46, 20, -79, -99, 40, -16, -1, -105, 104, 94, 122, 99, 8, -47, -125, -126, -28, -43, 45, 52, -114, 96, -63, 41, 87, 78, -118, -54, 124, 3, -13, 43, -105, 36, 72, 64, -107, -56, 87, 125, -90, 81, 96, 46, -94, 100, 48, 6, -71, -35, -70, -57, -66, -4, 112, -107, -54, 123, -32, -58, -2, 83, 113, 21, -8, 58, -43, 13, -126, -84, 10, -88, 126, -21, 86, -96, -49, 6, 39, 8, 100, 97, 80, -94, -35, 64, -73, 39, 59, 23, 110, -71, -21, 95, 79, 99, 25, -92, -16, 27, -47, 122, 67, -49, -27, 25, -17, 52, -96, -106, -67, -124, 120, -115, -90, -43, 77, -35, 125, 9, 117, 107, 66, -32, 74, 17, -61, -28, 54, 51, 127, -121, 45, 67, -42, -109, -36, 69, 71, -4, 92, -124, 0, 84, -111, 38, -87, 95, -124, -90, -24, 121, -111, -86, -39, 92, 60, 28, -64, -14, -49, -65, -7, 124, -126, 79, -113, -33, 20, 87, 91, -16, 91, -36, -60, 109, -126, -18, 76, -122, 20, -76, 127, 38, -34, -40, 2, -102, 116, 66, 12, -61, -127, -123, -64, -124, 84, -49, -29, -23, -90, -66, 89, -126, 26, -98, 111, 29, 12, 59, 35, -96, 111, 35, 70, -51, 123, -56, -24, 112, -118, 116, -77, -116, 122, -13, -112, 78, 67, -13, -73, 105, 49, -111, 107, -52, -81, 90, 105, 59, 21, 12, 91, 4, -81, 34, 82, -85, 106, -70, -101, 117, -82, -50, -127, -88, 66, -111, 119, 5, 4, -82, -18, -75, -65, -38, 1, -18, -76, -22, -87, 74, 119, -123, -50, -90, 39, -96, -47, 17, -38, -20, 6, 9, 59, 7, 49, -3, 24, 40, -126, -100, 87, -16, -46, -106, 74, 83, 5, 127, -66, 46, 73, -75, 51, -105, -37, -38, -72, 45, 108, 18, -103, -14, -101, 84, 122, 77, -47, 18, -11, -45, 47, -52, 68, -127, -29, 14, 84, 104, 13, -110, 22, -42, -57, -54, -18, 35, 36, 38, -48, 16, -72, -23, -125, -44, -66, 125, -95, 15, 15, 22, 99, -66, 99, 39, -65, -58, -75, -108, -82, 67, -90, 68, -103, -18, -114, 7, -111, 51, -83, -31, -61, -26, 74, -58, 58, -120, -61, 91, 24, 83, -15, -5, -111, -44, -94, -47, 26, -41, -27, 72, -102, 11, 13, -76, 121, 27, 59, -118, -50, 105, -21, 18, -49, -74, 88, -119, -66, -100, 100, 86, 111, -43, -47, -128, 42, -13, -47, -60, 75, 54, -115, 101, -62, 26, -103, -69, -75, 85, -58, 4, 62, 49, -106, -115, 103, 110, -106, -90, -118, 122, 124, 121, -49, -50, 122, 121, 65, -53, -66, 12, -126, -53, -14, -60, 101, 11, -1, -102, -32, 69, 30, -98, -9, 52, -85, -34, 35, -63, 4, 45, -69, 1, 39, 11, 79, 33, 4, 16, 108, 66, -99, 110, -115, 15, -78, 114, -102, 50, -115, -5, -9, 43, 25, 110, -32, 69, -51, -125, -122, 81, 48, -62, -46, -41, 77, -95, 120, -47, 50, 101, -108, 79, 83, -95, -34, -122, -108, -8, 56, -95, 115, -81, 76, 13, -98, -84, -46, -21, -81, -40, -68, 96, 26, 15, -73, -25, 48, -80, 57, -30, -107, 77, -79, 104, 110, 15, 110, -126, -120, 38, -93, 123, 86, 112, 8, 116, -100, 90, -33, -52, -77, 27, -84, 77, -86, -29, -75, 91, 19, 110, -67, 40, 59, -17, 17, 41, 126, -1, 44, -122, -90, 79, -126, 124, 63, 10, 112, 92, -27, -49, -88, 24, 106, -44, -27, -107, 55, 26, 112, -53, 8, -83, 115, -61, 28, 4, 109, 27, -124, 25, 33, -86, -24, 35, -90, -88, -82, -106, -124, 19, -27, -84, -85, -49, 0, 16, -28, -73, -85, -44, 2, 51, 2, -10, 119, -98, 122, 100, 57, 126, -3, -37, -88, 101, 126, -50, -115, -84, -28, -111, 63, 73, -67, 106, -103, 61, -5, -3, 117, 38, 82, -9, -39, -44, 109, -48, -14, 104, -76, -84, 102, 49, 7, -113, 23, 5, -35, 36, 50, 66, 54, -15, 11, 115, -36, 36, 49, 87, -94, 38, -3, 116, -99, 86, -56, -117, -89, 58, 115, -37, 102, 89, -115, -19, 104, 36, 115, -58, -56, 37, -120, 126, -106, 19, 114, -14, -72, 35, -55, -38, -55, 70, -50, -26, 29, 22, -15, 68, -48, -28, -97, -73, -66, -84, 36, -90, 80, 23, -20, -103, -68, -12, -105, -45, -120, -119, 69, -64, 44, -113, 26, 117, 85, 104, -36, -14, -2, 77, -74, 78, -78, -42, -123, -16, 2, 42, 22, -45, -63, -125, -20, -2, -9, 3, 81, -1, 13, 22, 63, -71, 37, -39, -81, -5, -63, 11, 109, 63, -40, -92, 14, 10, -6, 19, 122, 124, -67, 17, -49, -1, 20, 59, 125, -117, -65, 78, 11, 76, -28, -54, -123, -118, 36, -76, 5, 101, 63, -14, 37, -104, 22, -77, 34, -112, 70, 29, -115, -124, -82, -36, 3, 66, -104, 0, 77, -41, -50, -40, -93, 50, 35, -88, 60, -57, -35, -63, -84, -100, 52, 81, -76, -54, -124, 87, -37, 75, -12, -24, 79, 34, 68, -46, -28, 92, 82, -79, -77, -96, 10, -42, 82, -83, -1, 15, -12, 92, 80, 32, 120, 4, -14, -83, 79, -10, -124, -86, -63, -8, 18, -112, -102, -42, -30, -2, -77, -76, 47, -26, -44, -71, 61, -89, -26, -68, 54, 90, -104, 6, -5, -112, -117, 109, -67, 90, -29, -63, -124, 37, 57, 22, 53, 83, 108, -104, -47, -97, -52, -127, 6, 33, -70, -61, 72, 33, -1, -2, -5, 23, -124, 118, 39, -113, 99, 101, 105, -57, -90, 109, 108, 96, 3, 33, 51, -16, 57, -123, 15, -122, -122, -107, 39, -64, -40, -17, 97, 87, 109, -35, -18, 113, -45, -106, -127, -73, 123, 106, -2, -95, 88, -22, -127, -37, -117, 53, 75, 69, 58, -37, 75, 64, -16, -14, -128, 73, 97, 98, 32, 78, -65, -113, 63, 18, -91, 64, 73, -96, 43, -57, -63, 3, 49, -61, 94, 61, 120, 42, 2, 50, -123, -51, -14, -11, 63, -14, -66, 32, -44, 95, -18, 19, 110, -83, -90, -109, 110, 111, -77, 25, -73, -12, -100, 104, 55, 122, 37, 47, 36, -89, -31, 41, -12, 83, -97, -77, -58, -35, 83, 26, -68, -63, -82, -86, -17, -44, -67, -35, -61, -16, 118, -6, 101, -110, -29, 28, -116, -120, -52, 49, -80, 45, -38, 36, 1, -7, 88, 71, 87, 43, -31, -109, 109, 15, -66, -36, 99, -5, 57, -89, 108, 47, 33, 81, 65, -124, -19, 77, -115, 57, -2, -67, -25, 89, 97, 104, -46, 57, 47, -87, -27, -112, -67, -46, 32, -5, 46, 3, 118, -25, 42, 98, -106, -52, 51, 87, -48, -95, 36, -35, 90, -93, 26, -63, 124, -4, -87, -50, -75, 88, -8, 26, 105, 53, 108, 9, -80, 26, -116, -90, -127, 55, -119, -105, -125, 60, 110, -45, 93, 19, 49, 56, 54, -53, 121, 50, 71, -93, -128, 125, 123, -8, 23, 100, -83, 4, -19, -35, -98, -6, 4, -96, -79, 13, -73, -76, -55, -90, 7, -89, 57, -72, 95, -17, 4, 88, -95, -53, 123, -95, -56, 119, 26, 96, 91, 71, -28, -55, -91, 2, 67, 41, 34, 116, -74, 90, -88, -1, -128, 47, 38, 57, 104, 5, -88, -20, -34, -55, 55, -39, -22, -128, -48, -124, 96, -84, 76, -60, -11, 113, 70, -72, 26, -23, -84, 80, -61, -44, -49, -61, -125, 118, 124, 107, -5, -92, -41, 89, -19, -113, -77, 87, -113, 3, 92, 111, 47, 40, -77, -92, 25, 121, -36, -77, -30, 8, -125, 37, 92, -46, 104, 96, -56, 100, 75, 68, -120, -93, 29, -11, -78, 80, -51, -63, -44, -87, -80, -125, 81, -29, -88, -22, -36, 4, 29, 63, -115, 32, -28, 105, 114, -51, 73, -69, -79, 21, 127, -70, 56, 28, 47, 106, -19, 124, -85, 65, -91, -37, 68, 118, 62, 108, -32, -102, -15, 125, 89, -2, 29, -66, -25, 16, 11, -79, 75, 60, 70, 74, 118, -2, -26, 38, -24, 83, 34, 19, 20, 72, 110, -39, 62, 44, -59, -97, 70, 54, -100, 32, -76, 58, 94, 28, -54, -23, 77, -107, -91, 19, 95, -100, -111, -59, 66, -7, -103, -28, -116, 45, -84, 122, -122, 107, 38, -52, -118, -20, -126, -90, -116, -73, 96, 106, 83, -86, -45, 32, -65, -7, -77, -98, 21, -60, -28, -41, 61, -3, 59, 73, -86, 104, 67, -79, 83, -23, -3, 93, 85, -1, -125, 98, 54, 100, 76, 9, -114, -96, -87, -50, 25, -36, -20, -82, 32, 80, 5, -35, -51, -64, -90, -8, -88, 105, 41, 123, -46, -90, 88, -88, 37, 92, -118, -36, 64, 86, 101, 78, 118, -113, -100, 15, -21, 9, 61, -116, -39, -62, -23, 39, 3, 16, -97, 43, -7, 72, 39, 76, 110, -1, 116, 19, -37, 126, 111, -101, 84, 85, 106, 75, 100, -122, -38, -49, 15, -104, -37, 105, -38, 69, 16, 93, -43, 47, 9, 78, -9, -80, 26, -27, 47, 14, 120, -117, 12, 104, -90, -31, 61, -112, -84, 33, -105, 6, 112, 38, 30, -52, 15, 121, -111, -97, 86, -26, 78, -33, -76, -59, 15, 79, 42, -65, -35, 35, -54, 106, 11, -16, -53, -56, 1, -9, 105, 24, 125, 89, -66, 28, -91, 78, 21, -74, 109, -21, 28, 60, 75, 81, -127, -38, 32, 44, 25, 125, -49, 99, 103, 90, -44, -78, -94, 85, 41, -117, -19, 39, 100, 43, -61, -118, -7, 88, -64, -25, -61, 93, -93, -114, 46, -92, -23, -50, 80, -126, -53, -97, 102, -77, 121, -70, -27, -101, -113, -113, -90, -4, 54, -117, -89, 121, -107, 33, 81, -43, -120, -108, -78, -85, -93, 96, -49, 12, -82, -96, 14, -6, -65, -12, 45, -71, 46, -110, -44, 61, -95, -5, -71, 87, 6, -31, 80, 27, -126, 33, 112, -118, 54, -93, -75, 89, -125, 4, -27, -78, 36, 115, 44, 100, -24, -39, -99, -106, -21, -15, 84, 13, 108, -115, -28, -14, -18, -75, -115, -16, 86, 126, -6, 12, -95, 47, -27, -92, -76, 74, -42, 88, 62, -126, 60, -90, -37, 89, -68, 71, -53, -112, -44, -73, -98, 56, 42, 12, 109, 55, 125, 68, 53, -9, -48, 86, -89, 54, 123, -37, 0, -47, -77, -66, -44, 112, -28, 47, 73, 33, -10, -108, 49, 74, -52, 79, 3, 118, -36, -16, 45, -39, -76, -29, 80, 5, -71, 119, -69, -76, -46, 59, 6, 6, 122, 90, -10, -34, 9, -65, 127, -128, -44, 49, 74, 32, 0, -51, 22, 92, 62, -61, -75, 114, 38, -122, -9, 96, 125, 50, -108, -48, -18, 26, 86, -24, -12, -52, 70, 126, 11, 70, 126, 95, -9, 72, -1, 119, -106, -107, 84, 84, -39, -119, 70, 127, -113, -66, 95, -115, 112, 116, -35, -34, 14, -77, 70, -125, -1, 13, -127, -118, -45, 127, 106, 74, 71, -23, 65, 93, -1, 21, 49, 88, 31, -8, 87, 46, 54, 55, 59, 38, 43, -104, -123, -71, -53, 75, -68, 74, -40, -67, 85, 43, -68, 63, -11, -124, -88, -73, 97, 39, 76, 19, -1, -21, -117, -41, -102, 65, -114, 85, -25, 57, 110, -20, 114, -71, -72, -81, -124, 16, -20, 89, -68, 41, 24, 49, 45, 64, 104, 14, -24, 53, -95, 103, -96, -84, -66, -70, 109, -52, -112, -43, -123, 126, 65, 120, -73, 121, -89, -69, 10, 19, -108, 70, -68, 44, -9, 105, -19, -32, -8, 85, -107, 25, 60, -75, 70, 123, -16, 51, -57, 0, -120, -51, -2, 74, -59, 53, 67, -20, 113, -51, 127, -123, -109, -68, 50, 11, -91, -97, 107, 29, 116, -128, -73, 48, -75, 125, 43, 37, 48, 115, -91, 57, -64, 35, 3, 5, -39, -58, 113, -54, 20, 112, -49, 39, -84, -127, -78, -46, -96, -99, 111, -108, -99, -90, 69, -45, -93, -16, 120, 84, -29, -98, 13, 35, 65, -112, -88, -102, -42, -103, -28, 106, -118, 52, 18, -74, 53, 68, 8, 86, 98, -8, 106, 127, 30, 47, -46, 66, -96, -53, 22, 3, -23, -93, -89, -86, -77, -49, -59, 9, -23, 41, -12, -13, -35, -122, 41, -109, 74, -78, 105, 44, 42, 83, 44, -56, 3, 126, -118, 35, -55, 32, -90, 50, 67, -51, 93, 118, 29, -94, 0, -122, 75, 116, -7, -87, 122, -94, -68, 68, -44, -91, -15, 126, 120, -99, -57, -5, -101, -47, -98, -27, 114, -59, -105, 53, 18, 116, 44, -81, -106, -84, -75, 98, -96, 46, -117, -102, 81, -57, 94, -91, -20, -49, -92, -28, -20, -21, 96, 8, 60, 126, 109, 46, -61, -124, -28, 86, 121, -112, -123, -113, -68, -69, 113, -36, 105, 124, -10, 58, -61, -44, 96, 47, 36, -124, -108, -112, -17, 116, 24, -85, 114, 5, 90, -74, 10, -66, -116, 3, -50, -111, 18, 10, -52, 4, 102, -74, 0, -36, 112, 68, 48, 80, -13, -44, 84, 7, -27, -61, -5, 125, -17, -18, 3, -55, 36, -115, 7, 48, 16, 85, 65, -94, -33, -114, 38, -59, -60, -89, 33, -76, 107, -47, -123, -34, 38, 89, 102, -117, -99, -31, -120, 12, 79, 11, 85, -13, 24, -36, -93, -88, -79, 101, -53, 16, 115, 113, 85, -73, -104, -10, -21, -125, 71, -16, -30, -19, -54, -56, -8, -25, 41, 1, 115, -7, -116, 72, 108, 37, -92, -112, 77, -43, 117, -104, 101, 104, -118, 58, -97, -94, -80, 10, -90, 119, 123, 8, -27, -59, 80, 93, 44, -7, -34, 31, 114, -21, -25, 95, -112, 11, 111, 93, 96, 100, 118, 69, 76, -128, -1, 107, -94, 47, -11, -56, 38, -16, 80, -117, 53, 32, 105, -31, -102, -57, -128, -116, 50, -25, 107, 66, 114, 90, 32, 82, 62, 22, 23, 10, 22, -106, -11, 56, 69, 107, -127, -20, -37, 81, -9, -111, -14, -32, -14, 12, 40, -13, 24, -38, 90, 4, -99, 77, -34, 61, 31, -99, -45, -73, 39, 105, -51, -99, 33, -109, -120, 34, -1, -29, -12, 118, -12, 102, -41, 103, -14, 127, -38, -118, -39, -76, 14, -10, -127, 109, -77, 33, -118, 6, 88, 49, -17, -91, 78, -111, -72, 86, 51, 55, -70, -89, 46, 46, -115, -123, 21, -1, -124, 111, 10, -35, -92, -104, 84, -91, -123, -121, 70, -113, 14, 30, 65, 125, 68, 15, -114, 124, -26, 66, 52, 32, 105, -30, -50, 119, -25, 100, -10, -21, 83, -128, 72, 119, -103, 28, -99, -98, 36, 99, -82, -78, 2, 111, -81, -58, -2, -66, -62, 100, -128, 118, 4, 105, -40, 83, 96, 63, 55, -41, -86, 10, -41, 115, 2, -16, 15, 31, 15, -77, 2, 61, -27, -124, 44, 21, -54, -86, 83, 13, -113, 83, 3, 19, 60, 92, -26, 29, 27, -99, 116, 70, 40, -53, 57, -86, 60, -56, 73, -53, -4, -53, -120, 97, -48, 52, -10, 26, 94, -55, -89, 109, -100, 43, 1, 89, 7, 103, -10, -94, -123, -22, 104, 45, 53, 33, 87, -15, 106, 32, 60, -26, 107, 68, -57, -69, -8, 62, 86, -41, -121, 125, -60, -92, 40, 69, 125, -81, 45, -13, -46, 50, 93, -70, -33, 18, 92, -74, -124, 70, 86, 64, -84, 65, 5, -13, 125, 125, -79, 83, -44, -71, 80, 25, -35, -7, -34, -38, 40, -117, 77, 122, 61, 42, -75, -100, -68, -111, -46, -64, 87, -88, -127, -125, 106, 6, -10, 103, 3, 40, 58, 88, 97, 10, -15, -66, -125, 79, 24, 44, 91, -27, 38, 24, -113, 91, 53, -53, 108, -121, 12, 67, -80, 13, 70, -102, -109, -67, -127, 22, 101, 59, -18, 70, -59, 95, -124, -55, 47, 28, 117, 10, -127, 27, -94, -112, -9, 87, -37, -29, 95, 103, -89, -113, -12, 109, -87, 7, -86, -86, -98, -113, 101, 12, 85, -86, -20, 89, -13, -101, -11, -24, 37, -10, -124, 71, 6, -5, 31, 98, 94, -2, 73, -123, 13, -66, 115, 54, 69, -99, 96, 99, -83, 69, -16, -126, 111, 92, 92, -29, 119, -47, 75, 28, 72, 79, -29, -50, -54, -126, -80, -87, 0, 122, -82, -115, -72, -95, 67, 125, -65, 35, 97, -20, -24, -47, -18, -40, -83, -54, 59, -92, 28, 6, 64, -28, -42, -93, 50, 32, -90, 99, 73, 38, 93, 120, 52, -107, -103, -9, -110, -40, -101, 115, 68, 3, -60, -77, 91, -15, -3, 22, 21, -103, -99, -43, -3, -13, -7, -80, -109, 31, -109, 93, -59, 112, 85, 121, -123, 110, -15, -105, -57, 12, -117, -117, -113, -49, -66, 107, 65, 60, 1, -42, 85, 30, 44, -45, -111, -91, 3, -91, 68, 22, -126, -119, 6, 87, -125, 11, 69, -12, 34, -116, -128, 45, -104, -113, 125, -42, 122, 62, -110, -4, -108, 104, -102, 64, -69, -84, 101, 62, -47, 41, -44, -45, 51, 90, -86, 54, -27, 111, -86, -121, 124, -86, 53, -108, -71, 50, -22, -76, -16, -3, 48, 4, -27, 74, -59, 32, 118, -86, -34, -57, 84, 50, 26, 7, 12, 68, -67, 113, 52, -25, 120, 48, 17, 45, 68, 74, -33, -82, 126, 79, 43, 46, -44, -112, -7, 25, 48, -17, 67, -114, 55, 23, 64, -47, -98, -52, -106, -37, -67, 74, 66, -74, -6, -45, 99, -66, -98, -61, -20, -100, -110, -104, 75, -26, -88, -60, 127, 89, 51, 67, 103, -22, -38, 40, 60, -7, 116, 82, 84, -78, 28, 23, -24, -106, 106, -53, -44, -120, 14, 64, -91, 33, 88, 112, -121, -127, -76, -121, 90, 103, 74, 65, -46, -92, -23, -114, 29, -34, 96, -14, 16, -4, -119, 120, 18, 115, -61, 102, 124, 82, 38, -95, -13, -1, -111, -6, 0, -59, 1, -38, -84, -53, -101, -2, -16, 5, 12, -115, 99, -20, -1, -13, 104, 8, -21, -6, -4, 46, -32, -8, 0, -121, 25, 115, 6, 42, -18, -122, 111, 111, -32, -101, -69, -5, 26, 43, -128, -90, 56, 99, 19, -72, -42, -5, 64, 65, 118, -68, -16, -42, 52, 112, -35, -51, 100, 99, 119, -46, 105, 102, -63, -55, -126, -4, 69, 28, -89, 69, 66, 96, 41, -43, -104, 127, 81, 88, 65, 71, -107, -79, -99, 73, -95, -5, -105, -123, -34, -114, -41, -56, 117, 25, 17, 119, -107, -42, 19, -67, -100, -43, -99, 69, 43, -75, 68, -4, -115, 5, -61, -94, 54, -32, 108, 88, 91, -125, 93, -70, -111, -75, 2, -122, 78, -109, 125, 99, -22, 16, -96, 6, 102, -67, -53, 17, -14, -113, -115, 0, 21, -48, 34, -53, 48, 14, -93, 12, 17, -127, 70, 35, -74, -56, 41, -124, -37, 39, 103, 69, -73, -120, -53, -99, -59, 22, 46, 56, 38, 59, -72, -69, -117, 90, 6, 60, -23, 42, -56, 122, 43, -114, 29, 97, -42, -57, 101, 49, 110, 76, -9, -91, 84, 66, -61, -102, -39, 113, 82, 127, 45, -118, -70, 56, 100, 64, -12, -51, -22, 60, -56, -107, 74, 101, 118, -96, -84, 91, 82, -102, 40, -55, -64, -4, -117, 3, 22, -28, -12, -24, -29, -95, -14, 29, 90, -41, -34, -50, 36, 72, -117, 108, 94, 85, 82, 84, 118, 126, 48, 72, -103, -40, -111, -39, 84, -100, 92, -21, 1, -48, 83, 100, -14, -58, 2, -52, 29, 96, 26, -63, 40, 37, -82, 6, -5, -128, -37, -15, 126, -117, -71, -105, -29, -54, -16, -73, -26, -52, 34, 103, 29, -10, 76, -113, 60, -50, -37, -39, -82, 117, 26, 86, 27, 72, -35, -106, 72, 56, 7, 71, 67, 64, 94, -90, -118, -49, -35, -16, 27, -128, -40, -72, -10, -92, -57, -78, -14, 34, 11, 32, 24, -91, -10, -77, 110, 83, -55, 54, 11, 80, -3, -50, 16, -36, -12, 26, 43, 82, -118, -58, 82, -30, -1, -56, 6, 70, -6, 120, -23, -123, 24, -127, -86, -113, -76, -104, 98, -3, 79, -18, -51, -52, 60, 93, 40, -79, -9, -45, -125, 1, 26, 85, 100, -103, -99, -22, 95, 23, -29, -56, 28, 123, -55, 70, -118, -3, 95, 109, 122, 46, -37, -57, 122, -105, -92, 35, -56, 27, 118, -53, -99, 16, -96, -127, 41, -67, -21, 9, 84, 78, 81, -16, 74, -101, -73, 84, 24, -106, 65, 19, 68, -100, 90, 62, -76, 127, -31, -4, 26, -40, 72, 55, 104, 104, 56, 18, -90, -92, -101, 122, 114, 108, -21, 60, -121, 34, 17, 32, 56, -46, -77, -4, -17, -115, -70, 35, -116, 28, -97, 39, 116, 103, -34, 92, 80, -105, -18, 118, -69, 9, 112, -83, -10, -37, 106, -3, 125, -5, -99, 53, 77, -48, -79, -68, -34, -20, 95, -22, -120, 127, -111, 124, 102, -16, 88, 54, 7, -57, 44, 66, 80, 29, 111, -58, 120, 89, 68, 118, -44, 97, 43, -94, -78, 93, -34, 16, -55, -66, 122, -47, -67, -116, -51, -93, -4, -91, 90, -125, -20, 6, 69, -67, -93, 52, 3, -100, 14, -57, -110, 98, -87, 61, -124, -37, 26, -29, 107, 99, 33, 101, -76, 94, 113, 1, -127, -19, 39, 91, -16, -109, -30, -75, -48, 5, 106, 84, 33, -8, -101, 51, -38, -60, -15, -33, 31, -117, 66, 10, 111, -29, -16, -93, -63, -31, 37, -62, 79, -52, -98, -65, -33, 0, -11, 48, -123, -33, 4, 39, 87, 31, -38, -79, 100, 75, 16, 3, 87, -46, -114, 70, 53, -2, 105, 118, 95, 14, -71, 46, 90, -41, 110, -70, 87, -29, 106, 92, 66, -18, 3, 25, -115, 94, 74, 113, 41, -37, -11, 0, 45, 3, -58, -29, -127, -80, -39, 96, 62, 18, 15, 25, 105, -3, 83, 64, 96, 61, 29, 34, -85, -96, -69, -72, 126, -123, -86, 40, -32, 31, -88, -114, -94, -17, -15, -93, 31, 74, -125, -35, -35, 18, 118, -58, -113, 73, -121, 111, 6, 36, 17, 49, 68, 76, 106, 67, 82, -108, -21, -78, 51, 19, -64, 85, -126, 49, 120, 33, -4, 123, 127, 89, 14, 117, -97, 29, 63, -90, 13, -59, 74, -98, 119, 15, 107, 97, -46, 61, 117, 61, 111, 40, -48, -80, -3, -45, 97, -11, 116, -35, -16, 115, -74, 126, 105, -42, 28, 40, -4, -87, 109, -57, -57, 100, 86, -78, 69, -88, 111, 58, 101, 95, -30, -75, -113, 95, 8, 112, -44, -3, -50, 69, -16, 4, 67, -39, 90, -33, -127, -41, 8, 111, 30, 80, 83, -12, -126, 25, 28, 114, -45, 1, 81, 54, 54, 96, 21, -65, 80, 106, 60, -98, 47, -84, 35, -14, 6, -3, 82, 7, 84, -38, -10, -14, -86, -54, 102, -83, 99, 2, -97, -74, -125, 112, 108, 58, 80, 2, 121, 32, -20, 53, 63, -101, 97, -30, 13, -25, 95, -33, 111, 52, 58, -27, -90, 100, 47, -115, -111, 18, 15, -80, 73, 19, -96, 53, -51, 112, -73, -58, 17, 35, 123, -48, 62, 92, 50, -52, -60, 17, 43, -77, -59, -27, 24, -20, -54, -56, -7, -37, 90, -120, 12, 35, 27, 44, -39, 104, 29, 16, -82, -82, -76, -87, -2, 114, -122, -80, -66, -54, 65, 106, -3, -121, -49, -107, -13, 25, -35, 108, 117, -72, 116, 1, 91, 16, -83, -76, -8, 74, 69, 39, 120, 121, 80, -10, 107, 86, 38, -86, -96, -24, -108, 29, -17, -29, 51, 98, 125, -112, 78, 114, -56, 66, -13, -92, -46, 32, -40, 75, -21, -99, -14, -29, -106, -62, 90, -126, -103, 0, -84, -71, 104, -64, 87, -41, 35, 10, -71, 32, 26, -121, 18, 99, 74, -123, -121, -100, 38, -33, 103, -111, -3, -39, -12, 19, 28, -50, 21, 53, 79, 65, 110, 55, -127, 69, -113, 37, -49, -56, -59, 106, -48, 88, 77, -102, 93, 84, -74, 3, -77, -98, 20, 48, -9, -119, -60, -109, -41, 89, 72, -90, 27, 55, 94, 28, -4, 109, -63, 76, -75, 7, 54, 5, -33, 3, 31, -68, -41, 86, 64, 10, 116, -44, -69, -21, -35, -1, -1, 53, -40, -57, 91, 115, 126, 57, 16, -5, 38, 81, -57, 92, -40, 125, -31, 55, 0, -127, 116, 87, 87, 52, -31, 75, -120, 28, -74, -26, -101, 53, -101, -12, 125, 118, -25, 123, 48, 119, -10, -42, 73, 61, -78, -95, 58, 20, 89, -70, 21, 77, -111, -20, 1, -13, -73, 9, -113, -19, 111, -85, -93, -118, 31, -96, -127, -122, -101, 49, 126, 18, -121, 71, -49, -70, 104, -118, 78, 65, -60, -29, 14, -42, 79, -113, 73, -122, 25, 88, -13, 8, -125, 22, 19, 34, 54, 20, 41, 82, -59, 39, -28, -52, -18, 51, 6, -42, 61, -44, -104, -126, 55, 38, -40, 6, 54, -95, 12, -49, 121, -128, 87, 125, 22, -22, 31, -51, 126, -56, -97, -61, 111, 3, 16, -35, -74, -106, 52, 116, -21, 76, 118, -94, -14, -50, 41, -88, -17, -75, -9, -24, -75, -49, -27, 76, 57, -123, -103, 56, -51, -72, 123, -67, 59, 11, 26, 113, 34, -50, 101, -115, -102, 91, -81, 13, -87, 88, 53, 24, -114, -83, -127, -61, -4, -26, -113, -75, -21, -88, 109, 57, -32, 105, 118, -101, -12, 16, -115, -106, 95, 114, -93, 121, 78, -45, 6, 119, -85, -68, 16, -71, -23, 17, -3, 101, 119, 12, -102, -29, 53, -120, -100, -107, 113, -110, -79, -27, 34, -66, -4, 1, -80, 31, -5, 126, 114, -127, 118, -98, -67, 6, -41, 38, -105, 84, 11, -114, -31, 38, -15, -106, 46, 13, -85, 31, 31, -36, -124, -62, 26, 0, 67, 75, -96, -66, 73, -110, -64, 63, -80, -3, -59, 8, -92, -36, -36, 47, -21, 61, -43, 92, 83, -125, -22, 127, 34, -119, -37, 39, -53, 118, -89, -113, 65, -57, -51, 10, -38, 13, -54, 10, -117, 15, -110, -81, 108, -17, 94, -41, -84, -76, -77, -128, -73, 29, 127, 90, 39, -38, 1, 114, -48, 40, -127, -111, 112, -49, 28, -54, 92, 102, 84, 103, -11, 103, -106, -31, -42, 117, 56, 2, -87, 108, 2, -32, 9, 1, -70, -80, 92, 59, -93, -84, -28, -92, -66, -44, -13, 90, 30, -48, 64, -14, -73, -75, -39, -50, 23, 47, -61, -49, -78, -20, -69, 52, 76, 69, -74, -121, 117, -110, 66, -104, -66, -90, -67, -4, -6, 48, -42, -104, -128, -106, 11, -72, -52, 100, 6, 99, 20, 73, -78, 70, -75, -18, -6, -127, -77, 48, -120, -88, 66, 75, -63, -127, 113, -2, -3, -20, -82, 84, 4, -81, 106, -113, -25, -74, 116, 109, -103, 8, 54, -52, -50, 107, 58, 72, 108, 109, -7, 117, -107, -69, 64, -42, -68, 49, 84, 58, -99, -125, 14, 34, -78, -8, 49, 25, 47, 37, 6, 72, -83, -68, -108, -5, -89, 78, -60, -109, 59, 61, -120, 81, 120, 72, -89, -75, -6, 124, 111, 23, 127, -3, -71, -79, 117, 107, 74, 36, 16, -48, -19, 62, 12, 1, -71, 51, -48, -3, 70, -117, -70, 79, 92, -77, 23, -124, -24, -111, -128, -41, 41, 127, 84, 98, -80, 73, 77, 122, -18, -34, -54, 91, -100, 86, -36, -43, 9, 44, 83, -49, 56, -115, -98, 20, -64, 54, 24, 40, 71, 24, 127, -16, 23, 83, -45, 71, 29, -96, 65, -117, -2, -117, 102, 26, 97, -62, 112, -22, 111, 67, 58, 39, 80, 88, -69, -111, 14, 84, 57, -42, -20, 57, 70, -124, 12, -103, 75, -87, -70, 13, -76, 56, 24, -102, -45, -6, -35, -61, 100, -52, -122, 30, 115, 86, -9, -82, 103, -123, -126, 33, -37, -17, -38, -94, -13, 102, -69, -66, -112, -11, 75, -60, -82, -28, -33, 1, 94, 60, 68, 66, -120, 74, -31, 123, 32, 88, -87, 8, 93, -84, -87, -71, 27, 3, -37, -114, -23, 22, -52, -7, -116, -104, 62, -70, -4, -99, 59, -38, 89, -1, -100, 97, -55, -3, 92, 105, -43, -123, -15, -77, -79, 26, -20, 76, -99, 71, 90, 7, -35, -89, -128, -23, -65, 62, 35, 59, 91, -34, -107, 52, 93, -79, 21, -90, 47, -15, -112, -124, -9, 1, -73, 40, -100, 35, -11, -71, -22, -49, 64, 72, -10, 65, -79, 53, -1, 85, -16, -37, -77, 5, -113, -111, 55, 37, -73, -26, -106, -57, -22, 13, 73, 34, -74, 101, -59, 43, -98, 48, 122, 95, -8, -15, 32, 41, -90, -97, -2, 23, -6, 50, -100, 10, 67, 83, -81, 122, -71, -59, -62, 36, 83, -117, -58, -119, 112, 11, 52, -114, -69, 46, 109, 51, -97, 13, -35, -58, 45, 91, 93, -89, 13, 121, 49, -48, 77, 96, -53, -122, -90, 13, 42, 121, 24, 112, -126, 8, -4, 54, 22, 55, -28, 4, -21, 4, -111, 72, 74, 62, 35, 39, 102, -79, 32, 23, 1, -19, -8, 76, -12, 30, -39, -98, 23, 113, -113, 25, -7, 11, -49, -112, -62, 51, 20, 45, -73, 37, -11, -127, -28, -103, 40, -54, -54, -55, 97, 75, 54, -39, 24, -86, 119, 113, -55, 14, 99, -40, -89, -36, 99, -10, -20, -91, -86, -128, 83, -31, 38, -56, -29, -118, -31, -117, -44, 43, -44, -75, -9, -117, 15, -113, -75, 6, -128, -2, -107, 99, 86, -68, -64, 57, 51, 44, 95, 93, 45, 50, -66, -45, 122, 33, -35, -36, 45, 49, -121, -127, 102, -2, -116, -11, 13, -62, 124, 14, 64, -111, -15, 23, -51, 49, -48, -128, -34, -81, 93, -117, 97, -100, -34, 92, 61, 59, -72, -22, -20, -65, -20, -46, 62, -8, 72, -53, 58, 68, 89, -5, 85, -53, -110, -94, 124, -30, -93, -38, 18, -128, -27, -13, -100, 67, -49, 90, -2, 7, -60, 106, 71, 48, -67, 5, -87, -123, 80, 99, 73, 42, -34, 30, 117, -16, 64, 113, 83, 99, -52, -27, 100, 49, 88, -128, -11, -88, 90, 115, 47, -97, 94, -10, 79, -101, 123, 120, -96, 76, 92, 105, -10, -70, 7, -21, 43, -57, -36, -2, -85, 40, 99, -113, -38, 59, -113, 79, 99, 106, 66, 19, -119, 32, -119, 88, 59, -123, 81, 91, 81, 45, 68, -57, 103, -53, 50, 18, 19, -114, -112, 62, 55, 115, 77, -111, 47, 92, 96, 18, 70, 34, -91, 79, -61, -81, 40, 126, -76, -7, 90, -123, -90, 30, -52, -115, 106, 126, 32, -3, -116, 48, -69, 67, 36, -120, 84, -45, 100, 52, 101, 43, -41, -117, -6, 26, -70, -94, 24, -18, 27, -14, -13, 65, -111, 63, 79, 123, 61, -17, -8, 73, -97, 51, 13, 67, 59, -31, -106, 31, -106, 124, -54, -19, -121, 69, -121, -63, 103, 31, 47, 3, -110, -94, -60, -93, 97, -109, -98, 30, 2, 22, -25, 34, -55, 116, -27, -124, -42, -4, 35, -20, -8, 110, 89, -1, 51, 96, 64, 26, -1, -17, -99, 17, 17, -30, 52, -14, -11, 82, -112, 120, -24, -9, 26, 49, -20, 127, 53, 66, -5, -39, -82, 115, -57, -121, -14, 122, 103, -78, 20, -26, 33, 50, 120, -78, -108, 44, 36, 9, -1, 52, 1, 103, -84, -101, 25, 24, -101, -50, -38, 22, 39, 8, 10, 110, 15, 124, 104, -10, -81, -3, 92, 80, -81, 84, -125, -61, 1, 39, 76, -128, -36, -50, 103, 8, -23, 0, -96, 4, 79, -6, -101, -10, -126, 37, -27, 17, 33, -51, -121, 80, 74, 99, 33, 121, 56, 36, -68, -71, -53, -119, -71, 39, -41, -96, -81, 64, 33, -49, -59, -16, 73, -32, 102, 75, -123, -53, -36, 38, 25, -29, -9, -29, -57, -104, -35, 127, 60, 25, -72, -121, 34, -15, 47, 121, 17, 94, 58, -78, -82, 127, 34, 119, -33, 9, 67, -28, 84, -97, -118, -19, 3, 1, 81, 74, 25, -82, 73, -43, 71, -127, -35, -22, -14, -116, -29, -125, 106, -99, -74, -104, -100, 88, -112, -5, -31, 83, 95, -74, 114, 106, 35, -11, -21, -12, -65, -123, 34, -120, -38, -22, -119, 55, 84, -5, 67, -73, -1, 46, -43, 53, 70, -15, 13, 86, 109, 111, 41, 76, -91, 28, 54, 72, -111, -94, -67, -47, -89, 95, -39, 1, -55, -29, -71, -99, 94, 124, -43, -35, 42, 42, -110, -15, -101, 32, -57, -120, 15, 113, 85, 52, 13, 11, -4, 30, 45, 57, 111, 84, 25, -55, -42, 98, 44, 15, -128, 10, 11, -43, 104, -74, 127, 122, 39, -102, 26, 110, -93, -87, 95, 120, 93, -20, 3, -38, -117, -79, -109, 122, -123, 44, -61, -37, 15, 111, 106, 15, -6, -10, 100, -30, 44, 99, -36, -45, 125, 119, -63, -96, -96, -95, -104, 126, 13, 28, -40, 24, 77, -21, 19, 82, -104, 86, -82, 39, 70, -104, -74, -64, 14, -102, 34, -70, 125, 126, 13, 122, 117, 79, -101, -106, 112, -77, -108, -3, 79, -20, -106, 28, 87, 41, -17, 111, -1, 29, 22, -59, 53, 76, 5, -60, 102, -89, -2, 99, -90, -116, 94, -101, 91, 121, -79, 75, -84, -59, -56, 124, 49, -34, 24, 9, -121, -121, -8, 7, 36, -113, 76, -38, 91, -46, 30, 66, -7, -100, 37, 31, -88, 3, 59, -125, -4, 108, 78, 41, -78, -105, 37, 99, -11, -67, -20, -3, -59, 101, -124, 105, 116, 80, -61, 79, -94, 97, 17, 28, 126, -73, -69, -90, 58, 118, -86, -73, 99, 120, 96, -107, -113, 5, 120, 5, 66, -27, -126, -121, -54, -122, 113, -66, 86, -76, -115, 121, -106, 31, 21, -108, 86, 80, -70, 16, 71, -28, 71, 42, -35, 39, 63, -20, -84, 55, 113, 111, -100, 115, 118, -26, 121, 103, 36, 80, -100, 50, 73, -78, -47, -34, -58, -89, -82, 0, 55, 117, 101, -1, 31, -62, -90, -34, 46, -45, -106, 32, -62, -78, 19, -72, 25, 13, -96, -67, -35, -68, 111, -90, -18, -64, 4, 52, -25, 50, -76, -97, 40, -103, 30, -57, -37, 68, 38, -118, -105, 60, 42, -39, 110, -67, 18, 7, 74, 50, 69, -89, 110, 52, -51, -36, 117, 81, -112, -36, 4, -60, -5, -84, -34, -103, -13, 57, 94, -103, 67, 117, 85, -19, -49, 68, 43, 97, -53, -11, 19, -112, 29, 1, 69, 106, 93, 58, 60, 109, -106, -64, -79, 18, -20, 15, 43, 95, -55, 9, 121, -116, -1, 78, -6, 78, 18, -91, 47, 94, 26, -62, 110, -73, 67, 51, -94, 32, -19, 94, 13, 4, -98, 62, -106, 10, -50, 65, -23, 23, -53, -30, 35, 74, -79, -99, 24, 67, -62, -57, 33, 93, 9, 16, -108, -52, -61, -74, 108, 49, -108, -7, -75, -78, -73, -53, 60, 5, -116, -90, -100, -41, 8, 64, -95, 57, 93, 57, -3, -96, -128, -98, 125, 9, 46, -111, 85, 114, -56, 65, 35, -36, -70, 88, 15, -14, -93, -53, 119, -81, -15, -108, 7, 122, 84, 40, 51, 49, -30, -80, 81, -30, -49, 78, 108, 125, 96, 65, 111, -88, 3, 18, 4, 61, -22, -109, -81, 13, -33, -89, 61, 80, -69, -60, 74, -113, 108, -2, 64, -50, 46, 18, 49, 125, -32, 29, 123, -64, -34, 106, -24, 97, -3, 109, 31, 103, -128, 78, -11, -33, 117, -78, -80, -80, -10, 122, -65, -30, -8, -128, 49, -89, 18, -30, -92, 114, 127, -97, -77, -35, -118, 27, -65, 7, 8, 94, -18, 9, 44, 99, 104, 34, -107, -104, 82, 11, -109, -110, 110, 11, -110, 31, 50, 36, -127, 87, 22, -128, 118, 73, -35, -128, -27, 28, 7, 109, -6, 118, -10, -89, 89, -33, 73, 111, -9, 27, -6, 10, 45, -24, -106, 63, -121, 72, -29, -120, 31, 122, -120, 22, 67, -26, 22, -88, -126, -98, -106, -3, -108, 12, 36, 109, 107, -19, 92, -29, -120, -41, 109, 54, 63, -125, -11, 71, 76, 89, 79, -21, 83, 88, -127, 22, -66, 24, 63, -64, 54, 85, 61, 74, -31, -31, 55, -51, 78, 20, 48, 87, 107, 29, 13, 42, 33, -126, -15, -19, 91, -63, 88, 46, -103, 90, -59, -41, -14, -124, 23, -88, 89, -43, 114, -70, 54, 41, 7, 5, -67, -73, -36, -88, 85, 105, 83, -10, 107, -60, 99, 71, 5, 59, -11, 30, 21, 58, 117, -121, 62, 13, -81, 23, 98, -95, 82, 24, 75, -39, -99, -120, 17, -7, -79, -26, -30, -124, 92, -50, -56, 63, -107, 78, -6, 10, -20, -112, -59, -30, -105, -125, 111, -57, 27, 81, -24, -19, -23, -77, 70, 7, -68, -41, -128, -19, 61, -29, -15, 25, 49, 57, -40, 70, 7, 83, -48, 116, 99, 21, -42, 122, 25, -59, -63, -76, -106, 42, 33, -1, 93, -25, -122, -103, 63, -121, 6, -4, -22, 119, -106, -101, 49, -18, 97, -72, -63, -79, -84, -92, 71, 2, -97, -32, 71, -32, 20, 93, -118, -75, -35, 104, 28, -29, -127, -37, -22, 8, 88, 84, -1, 110, 111, -80, -36, 80, -23, 30, -126, 21, 66, 73, -104, 97, -87, 95, -62, 61, 61, -52, 114, -102, -76, 14, -3, -74, 106, 104, 62, 66, 60, -67, 48, 44, -18, -116, -4, 87, 42, -2, -20, -19, -57, 4, -50, -16, -28, 16, -83, -95, 93, -97, -69, -111, 46, 56, -57, 24, 32, -123, -38, -35, -61, -118, -119, 49, -106, 5, 8, 65, -124, 116, -82, -53, -7, -4, 60, 93, -115, 105, 126, 106, -119, -71, 123, 55, 113, -61, -49, 18, -56, 41, 111, 11, 51, 120, -68, 73, -3, 68, 10, 1, 57, 56, 77, -78, -75, 9, -113, -62, -14, -115, -84, -5, -58, -89, -78, -73, -22, 1, 73, 51, -86, 56, -66, 93, 48, -5, 39, -82, -65, -79, 47, 120, 106, -4, -86, -97, -123, -71, -31, -8, -58, 13, 115, 12, 52, -90, 68, -97, 39, 13, 82, 82, -58, -112, 47, 118, 11, -42, -92, 75, 8, 84, 67, -14, -48, 110, 17, -42, -89, 114, 78, -18, -1, 65, 122, -77, 103, 62, -46, 15, -52, -92, -31, 18, -75, -112, 8, 64, -25, 45, 11, 111, 1, -49, -31, 81, -67, 114, -89, -28, 100, 117, 82, -29, 55, 77, 22, 30, 11, 105, -83, 87, -115, 14, -23, -62, 31, 114, -125, -122, 31, 14, 117, -96, 93, -42, 113, -102, -56, -103, -1, -84, -114, -47, 15, 69, -98, -91, -28, 42, -114, 17, 1, -100, -96, 107, -34, 63, 93, -31, 69, -4, 112, 58, 28, 77, -112, 13, 104, -40, 38, -25, 4, 53, 56, -109, -6, 87, -72, 94, 1, -57, -16, -126, -29, 16, 109, 65, -49, 74, -93, -108, -58, -109, 78, 98, 96, 94, -16, 72, -74, -106, -81, 58, 75, 104, 77, -58, 63, -123, -92, -64, -52, 20, -62, 47, -92, -80, -15, -13, 122, 20, 7, -63, 39, -43, -93, 7, -77, 19, -48, -23, 42, -1, -93, -11, -25, 112, 59, -90, 118, 96, -26, -62, -12, 41, 114, 25, 89, -29, -116, 83, 119, 20, -108, 30, 105, -72, -91, -99, 75, -11, 6, -11, 117, 42, 107, -36, 26, 38, 3, 16, 6, 105, 83, 123, 18, 69, 20, -21, -88, 32, -65, -97, -76, -45, 61, -98, 11, 98, -69, -41, -40, 65, 76, -51, -21, 55, 41, -122, -34, -84, 22, 100, -106, -23, 95, 40, -82, -13, -108, -42, -108, -45, -11, -56, 38, -78, -26, -78, -107, 33, 9, -19, -29, -43, 58, 78, -115, -29, 84, -21, 16, -21, -49, 38, 84, -81, -50, -125, 34, -30, -39, 54, 53, 79, 127, -36, -127, -27, 14, -106, -121, -105, 3, -22, -20, -67, -72, -7, 33, -115, 100, -79, -8, -76, 87, -52, -29, -91, -49, -123, 8, 41, 60, -67, -8, 59, 25, -7, -96, -89, 16, -89, -66, -109, 17, 43, -47, 74, -92, 114, 87, -119, -93, -49, -67, 122, 27, 32, -97, 107, 37, 39, 20, -31, 101, -116, -100, -2, 5, -67, 38, -107, -28, 100, -87, 118, 15, -6, 64, 52, -20, 23, 61, 15, 102, 122, 9, 1, 26, 40, -20, -65, -48, -128, 33, -75, -116, 61, 51, 18, 122, -39, 39, -33, -66, 80, -43, 77, -54, -107, 1, 54, 44, -66, -59, 18, -72, 78, -109, 82, -9, 0, -110, 71, 0, 51, 124, 13, -16, 47, -97, -21, -119, 70, 74, -57, 23, -97, -108, 97, -76, 22, 24, 96, 84, 93, -14, -115, 44, 5, 95, -93, -123, 113, 106, 6, 36, 102, -109, -107, 21, -78, 0, 30, 120, -54, 101, 15, -23, 122, -15, 29, 16, -119, -3, -28, 102, 111, -15, 18, -12, -47, 53, -6, -62, 31, -128, 103, 5, -109, 124, -101, -59, -4, 57, -67, 70, 31, 77, -81, 25, -66, 76, -87, -57, -55, 13, -83, -72, 127, 64, 44, -48, -11, -90, 18, -107, -90, -7, 26, -71, -11, 53, -2, 113, -17, 60, 55, -114, 9, 102, 39, 71, 50, 80, -114, 123, -35, -69, -77, -36, 123, 96, 44, -15, -122, -65, 6, -83, 56, -96, -26, -82, 86, 101, -97, -59, 33, 87, -45, -86, 61, 122, 113, -16, 74, 127, -21, -89, -70, 31, 4, -74, -1, -80, 39, 5, -17, -83, 50, -88, -51, -103, -42, -93, 126, -11, -24, 31, -52, 59, 73, -118, 53, 58, -6, -1, 57, 101, 39, 115, 4, -85, -87, -125, -37, 80, 9, 75, 125, -69, 115, -53, -44, -55, -18, -46, 62, 87, 113, -117, 18, 58, -107, -56, -12, 15, 71, -83, -12, -18, -95, 121, 25, -54, 124, 117, -101, 5, 64, -104, 65, 51, -29, -107, 124, 82, -24, 58, 41, -39, 69, -69, -108, 90, 3, 8, -23, -53, 54, 94, 57, 87, 87, -45, -95, 83, -56, -68, -39, -120, -43, -102, 59, 56, -81, 55, 10, 23, -15, -77, 113, -73, -17, -123, -111, 114, 13, -5, -67, -61, -39, 119, -102, -80, -54, -68, -125, 18, -8, -36, 26, 77, -10, -43, 6, 38, -116, -112, -67, -3, -60, -82, 52, 51, -77, 70, 37, 65, -63, 99, -124, 26, 90, -97, 74, -92, -37, 77, 54, 83, -86, -48, 33, 32, 37, -89, -58, 49, -73, 4, -82, -5, 50, 99, -82, 102, 41, 84, 39, 106, 55, 43, 4, 17, 74, -50, 53, -91, -101, -21, 121, -59, 59, 26, 102, -32, 65, -84, -111, 120, 48, -65, -12, -29, -94, 34, -55, 75, -10, 112, 53, -83, 27, -71, 62, -26, 7, -13, 11, 35, 94, 4, 104, 25, -98, 78, 121, 95, 123, -118, 88, 43, -54, -52, -114, -20, 110, -41, -72, -27, -57, 109, 18, 99, -89, -47, -55, 46, 68, 84, -47, 35, -39, -70, -68, -9, -120, -74, -41, -125, -64, -81, 47, 10, -5, 61, 119, -23, -107, -81, 78, -36, -100, -31, -65, -61, 50, 8, 114, -10, -35, -61, -103, 54, -3, -42, -83, 6, 12, 4, 9, 76, 51, -72, -41, -82, 118, -50, 24, -117, -3, -26, -25, 25, 71, 39, 93, -7, -81, 79, 112, 12, -110, -119, -62, 16, -33, -16, -106, 107, 116, 31, 56, 40, 88, -113, 86, 78, -35, -18, 89, 90, 85, -64, -13, 28, 103, -48, -106, -105, -97, -122, 35, -78, -113, 102, 66, -17, -42, 88, -38, -54, -9, -110, 114, -49, -95, 73, -99, -2, -73, 118, -40, -116, -73, 76, 41, -98, -100, 63, -75, -68, 69, 89, -18, 84, 63, -80, -61, -107, -120, 30, -33, -1, 48, -46, 79, 82, -101, 108, -48, -46, 99, 41, -33, -102, -11, -120, -72, 17, 71, -18, 77, 12, -57, -69, -32, -122, -21, 36, -101, -13, -62, -6, 115, 114, 76, 66, 68, 103, 46, -107, -70, 17, 62, 25, 43, -77, 33, 100, 68, -24, -46, 18, 116, 25, 77, -44, 31, -71, 120, 58, 44, -70, -76, 31, -83, -127, -31, 113, 104, -112, -122, -94, 33, 68, 59, -51, 119, -36, -79, 60, 68, 3, -50, 56, -100, -101, -115, 59, -44, -123, -11, -127, -64, 41, 32, -19, 42, -126, -34, 19, -110, -27, 53, 51, -87, -15, -128, -95, 77, -79, 93, 18, 52, -85, -54, 80, -58, -41, 11, 27, -35, -128, 28, 29, 42, -68, -118, -44, -66, -24, 103, -48, 77, 29, -124, 119, -114, -124, -104, 91, -74, 117, -19, 106, -96, 56, 59, -26, -113, -58, -127, -20, -57, 29, -119, 113, 90, -109, -59, -104, -4, -83, -23, -55, 74, -19, -64, 88, -15, -40, 51, 39, -51, -95, 18, -19, 89, -51, 84, 104, 19, 85, -43, 90, -13, -34, 75, -51, -14, -111, -27, 110, -66, 78, -73, -120, -69, -8, 96, 45, 80, 19, -44, -98, 52, 102, 11, 13, -77, -33, -10, 71, -75, 75, 33, 40, -87, -19, 117, 27, -2, -38, 9, 60, -87, 65, 68, -28, -71, 36, -111, -119, -73, -26, -89, 108, -52, 51, -7, 0, -110, 111, -57, -57, 58, 104, 111, 100, -43, 100, -1, 83, -65, -119, 15, -24, 74, -45, 76, -125, 119, 94, -116, -81, -60, -76, -101, 16, 103, 20, -112, 121, 4, -41, -63, -66, -64, -80, -94, 21, -107, 34, -23, -44, 43, 120, 60, -11, -52, 8, -8, -61, -26, 4, -14, 42, 56, 13, -69, 31, -94, -53, 25, 38, 35, 90, 100, 99, -118, -121, -8, -97, 41, 97, -13, -44, 90, -81, 73, -90, 56, -63, -23, -98, 69, 92, 73, -2, -23, -124, -99, 11, -49, 54, -79, 114, 16, -106, 85, 27, -99, -50, 58, 70, -81, -82, -102, -119, -35, 99, -81, -107, -92, 25, -76, 105, -11, 125, -25, 94, -127, 5, -22, -48, -69, 27, -61, 76, 49, -104, -25, 78, -26, -95, 20, 22, -49, 46, 31, 45, 17, 79, 66, 53, -24, 118, 31, 93, 115, -122, 59, 116, 11, -91, -59, 71, 65, 8, 19, -14, 32, 122, -63, -121, -101, 85, 29, -21, 4, -68, -104, -107, -117, 90, 75, -13, 81, -22, -48, 68, -16, -116, 57, 124, -79, 126, 67, 114, 6, -42, -27, -90, -48, 38, -83, -21, -5, 74, 86, 127, -121, 110, -107, -110, 73, 96, 6, 26, -54, 86, -34, 58, 98, -105, 54, -108, -107, -7, -122, 27, 79, -21, 66, -97, -111, 111, 11, 13, 58, -31, 12, 65, -48, 33, 83, -103, 1, -39, 51, 75, -80, -111, 6, -110, -87, -68, -90, -66, 54, -83, 90, 5, 24, 28, 37, 42, 11, -80, -73, -59, 17, 67, -122, 97, -27, 90, 122, 102, -77, 45, 50, -29, 63, -72, -10, 104, -12, 28, -90, -86, 73, -128, 48, -30, 28, -43, -116, -88, 5, -61, -19, -106, -122, -12, 120, -21, -50, 114, -46, 1, 32, -124, 101, -33, -68, -37, -57, 48, 119, -19, 91, 65, -18, 11, -93, -118, 96, -81, -78, -27, -14, 32, -5, -8, -108, -13, 100, -30, -26, -74, 99, -122, -70, 72, -27, -10, -93, 44, -90, -101, -103, -127, 92, 7, 12, 127, 18, -20, -82, 68, 81, 32, -28, -51, -104, -8, 64, 124, 90, -90, -78, 62, -84, -20, 6, 17, 98, 42, -67, -119, 69, -41, -118, 33, 94, 23, 32, -16, -125, 78, -75, 85, -18, 25, -94, 6, -110, 98, 3, 108, -119, 53, 42, -75, -94, -79, 71, -124, 91, -124, -115, 32, -37, -104, -63, -70, 47, 97, 42, 50, 47, 95, 7, -99, -7, 41, 35, 11, 12, -90, -9, 21, 92, -94, 74, 126, -45, 17, -126, -82, 22, -112, 78, 113, -88, -113, -85, 87, 112, 86, 9, 31, 53, -111, 60, -82, 58, -33, 57, -58, 6, -79, 91, -30, -45, 38, -32, 38, -73, -30, 84, 77, -14, 34, 63, 26, 49, 106, -15, 33, 64, 123, -64, -10, -116, 124, 36, 70, -37, -34, -115, 97, 15, 104, -61, 98, 14, 35, 8, 70, -122, -36, 19, -8, 126, -46, -109, 47, -67, 4, -48, 125, -1, 16, -13, 11, 12, -104, -46, 103, -10, -33, 73, -123, -57, -116, 103, 86, 48, -17, 28, 54, 75, -81, -82, 73, 2, -63, -8, 63, 70, 72, 60, -59, -40, -80, 81, 100, -56, -93, 75, 62, 2, 20, 67, 73, 33, 42, 31, -47, -103, -69, -121, 100, -21, -75, 45, 109, -9, -91, 44, -67, 109, -24, 2, -59, 24, -45, -87, 96, -10, 116, 30, 120, 9, -31, 66, -86, -117, -31, -5, -92, 29, 2, -120, -120, 55, 53, 117, -82, 90, 33, -21, 71, -119, 110, -116, 34, -63, -75, 2, 56, -86, -95, 48, 51, 2, -14, 93, 14, 84, -40, 50, -15, 90, 59, -7, 17, -16, -18, 64, -53, -113, -85, -110, -104, -103, -97, 58, -37, -44, -67, -109, -2, -34, 67, -79, 96, -74, -114, -18, -118, -26, -95, -5, -64, 92, 116, 82, -52, -30, 18, 23, -15, 61, 42, 9, 87, 73, -60, -78, -99, 1, -59, 28, 95, -120, 77, 63, -66, 92, -82, -56, -62, -49, 67, 3, -85, 55, -43, -9, -103, 103, -113, 10, 36, 57, -108, -5, 2, -40, 45, 31, 89, 114, -69, 56, 123, -119, -9, -71, 101, 37, 2, -89, 116, -59, 42, -97, 125, 127, 23, -106, 102, 38, 33, 11, -33, 53, -122, 97, -115, 52, 0, 102, 38, 60, 30, 33, 69, -107, 91, 42, 59, -35, 81, 47, 34, -4, 79, 31, -5, -26, 54, -30, -116, -41, 109, -21, -116, 115, -52, -103, 39, 76, 127, -50, 8, 29, 111, -51, 50, 74, 119, -19, -89, 73, -99, 74, -59, 108, -23, 64, -46, -97, -94, -34, -10, -113, 73, 2, -125, -107, 27, 42, 97, 26, 120, -22, -73, 104, 55, 106, 50, 47, -41, 90, -8, -12, 36, 61, -32, -115, -3, 50, -83, 32, -112, 35, 47, 89, -90, 50, 110, 65, -35, 80, -36, -43, -70, 19, -67, 113, -3, 112, 32, 85, 74, -104, -55, -18, 85, 42, -5, -45, -36, 40, 115, -19, -52, 34, -58, -14, -43, -75, -77, 50, -123, 15, -121, -65, -93, -59, -80, 32, -75, 81, -11, 127, 105, 63, -19, 63, -23, 104, -110, 69, 17, -123, -78, 93, 39, -7, -49, 124, 46, 2, 46, 51, -110, 54, 114, -75, 123, -94, 85, -80, 115, -53, -81, 93, -118, 28, 28, -13, 4, 46, -72, -107, 51, -21, 114, -38, 100, -63, -41, 18, 68, -123, -59, 86, 59, -73, -117, 54, -39, 96, 102, -51, -85, -107, -86, -75, 49, 70, 40, -74, -12, 97, -53, -89, -52, -66, 1, -80, -1, 88, 66, -61, 94, -121, -103, 25, -66, -92, -48, 23, -123, -74, 100, -80, -52, -114, -26, 125, 84, -114, -77, -56, 111, -1, -17, -69, 61, 113, -21, -68, 73, -83, 0, 39, -76, 25, -63, -14, 62, 17, -118, 67, 71, 110, 115, -109, 125, -39, -111, 81, -24, -60, -102, -41, 67, 9, 19, 0, -6, 126, 61, -60, -84, -67, 107, -32, 86, -84, 83, 20, 61, 93, -41, 5, 75, -53, 24, 72, 36, 41, 26, -116, 110, 52, -28, 49, -67, 119, -78, 56, 117, 111, 124, -95, -84, 103, 2, -126, -108, -43, 23, 81, -78, 110, -42, 125, -71, 111, 70, 94, 24, -32, 106, 6, -108, -50, -72, -47, -59, -22, -119, -69, -39, -123, -36, 5, 109, 94, 7, -127, -77, -98, 82, -27, -115, -87, -29, -58, -104, -87, -92, 48, 9, -113, -73, 29, -35, -17, 110, 35, 89, 120, 94, -78, 125, -70, 55, 106, -103, -66, 107, -52, -35, 62, 50, -22, 103, -107, 48, 127, -66, 85, 47, 71, 100, 102, -28, -63, -43, -46, 100, -82, -54, 66, -32, -56, 125, -105, -78, -106, -42, -98, -30, 51, 92, -108, -99, 67, -87, 77, 66, -25, 34, -15, -82, 6, -40, 18, 72, 45, 101, 44, 92, -81, -17, -68, -9, -20, -44, 42, 2, 42, 72, 100, -35, 36, 121, -6, -25, -94, -57, -87, 10, 106, 26, 56, -16, 114, -53, -72, 32, -80, 101, -4, -33, -44, 56, 87, 64, -116, 1, -62, 54, -55, -90, -109, 109, -97, 13, -44, -62, 85, -3, 76, 63, -105, 4, -81, -118, 79, -24, 42, 127, -51, -90, -33, 33, 94, -74, -31, 107, 55, 35, 33, -128, 73, 53, 109, 105, -62, -63, -85, -105, 62, 119, 86, 85, -5, -122, 95, -53, -18, 9, -54, 59, 47, 41, -36, 14, 95, 61, -7, 22, -32, -102, 22, -87, 79, 3, -110, -110, 68, -67, -87, 2, -76, -128, -40, 48, -122, -73, 123, -12, 65, -59, -81, -16, 111, 11, 126, 78, -56, -9, -27, 40, 18, 123, 81, -31, -1, 100, -13, -61, -95, 29, 70, -42, 29, -98, -122, 35, -43, -127, -105, -106, -58, -58, 7, -75, 81, 5, -124, -103, 125, -23, 65, 15, -28, 18, 112, 99, -10, -28, -89, 24, -127, 109, 110, 30, -117, 116, -63, -32, 117, -40, -9, -69, 30, 126, -15, -17, 3, -11, 8, 0, 94, -55, -113, -62, 91, -128, -90, -46, -28, -51, 106, -27, -70, 88, -125, -59, 76, -60, 37, 65, 28, -100, 124, -70, -102, -19, 41, 30, 98, -79, -98, 64, -6, -82, -125, -43, -82, -87, 39, 18, -10, 17, 119, 48, -23, 122, 117, -75, -66, 26, 118, 90, 55, 115, -108, 81, -32, 61, -17, -61, 110, 14, -125, -24, 60, -122, 61, 106, -81, -27, -4, 37, 118, -13, -43, -32, -19, -54, 21, 43, 101, 12, 5, 28, -1, 25, -19, 95, -42, 93, -94, -60, -21, -90, 44, -89, -84, -23, -111, -36, 78, 13, -127, 69, -128, -41, -91, -19, 33, 58, -104, 6, -58, 29, -94, 69, -74, 16, 37, 12, -19, 71, 80, 88, 109, -4, 127, -102, 101, -112, -10, 52, 29, -9, -7, 29, 78, 30, -118, -16, -40, -94, 118, 31, 63, -103, -28, 117, 41, -119, 1, -106, 81, -47, 110, 62, 77, 109, 88, 50, 125, -50, -26, 26, 70, 95, -73, 20, -3, -63, -124, 86, -29, 123, -11, -94, -108, 89, -105, 61, 99, 24, 83, 52, 105, 65, -14, 54, 46, -53, -24, 43, 25, 79, -59, -33, 46, -4, 116, -84, 61, 120, -126, -96, 115, -9, -62, -121, -48, -39, 68, -77, 113, 23, 103, 90, -40, -38, 16, -122, 37, 120, 49, -66, 71, 118, 30, -10, -14, 18, 34, -81, 10, 36, -49, -2, -101, 17, 5, -21, 106, -54, 31, 91, 97, 6, 53, -70, 96, -59, -64, 5, -66, 114, 68, -123, 104, -30, -5, -37, 116, -99, 10, -2, 65, 90, 124, 92, -21, 2, -56, -42, 76, 103, -79, 45, -19, 103, 103, -50, -84, -88, 83, -22, -102, 23, -16, -126, 121, 107, -35, 109, -119, 104, -20, 74, 66, -24, 39, -83, 106, 111, 3, 54, 86, 53, -28, -61, 28, -53, 17, 72, -13, -27, -77, 13, 124, 35, 16, 118, 14, 109, 99, 23, 85, -49, -30, 23, 56, -119, 69, 34, 120, -56, -39, 78, 125, 61, -111, 25, -120, 35, -30, -4, -120, 21, -119, -124, -72, 25, 122, 70, 7, 94, -34, -36, -83, 64, 116, 101, 73, 57, 8, 65, -127, 97, 15, 127, 30, 32, 24, 38, -61, 122, -94, -53, 15, -84, -48, 71, 69, -54, 14, -52, -88, 108, 41, -42, 44, 29, -69, -11, -42, 67, -74, -41, 36, 69, -42, -62, -27, 111, 105, 41, 105, -117, 116, -7, -73, -60, -64, 125, 15, 78, -55, 55, 58, 114, -115, -26, 15, -55, 91, 101, -116, -111, -67, 49, 86, 19, 115, -68, 2, 92, 101, -20, 104, 89, 101, -97, -98, -91, -100, 45, 116, -26, -28, 46, -40, -14, -107, 104, 59, 112, 77, 71, -126, -118, -8, 88, 30, -20, -108, -96, -56, 121, 12, -80, 83, -15, -48, 113, 23, -20, 30, 11, 82, -126, -71, -85, -12, -50, -109, -81, -65, 96, 119, -63, 107, -17, -103, 9, 91, -82, 41, -92, -89, -74, -44, 122, 39, 36, 107, -66, -111, 9, 73, 99, 12, -125, -114, -128, -47, -95, -80, 16, -126, -89, 81, 109, 22, 107, -10, -14, -103, -97, 22, -64, -43, 106, -69, 125, 15, -90, -69, 32, 48, -123, 3, -68, -120, 18, -68, -39, 51, -20, 106, 53, 19, 59, 34, -86, 38, -104, 28, 63, -72, -78, -128, 13, -100, -69, 10, 43, -31, 70, -53, -111, 75, 79, -51, 83, -31, 10, -84, -108, 118, -106, 74, 10, 82, -20, 52, -8, 5, -48, -72, 61, 2, -72, -54, 30, -13, 85, -54, 84, 27, 21, 102, -26, -28, -77, -71, 69, 61, -27, 90, 52, -4, 36, -66, -50, -112, 114, 70, 21, -62, 126, -46, 68, -74, 29, -30, 41, -14, 44, -2, -115, -62, -28, -13, 38, 23, 44, -20, -43, -111, -58, -119, 13, 106, -57, 91, 122, -71, 34, 16, -5, 32, 98, -65, 87, -1, 33, 0, 113, -50, 126, 126, 16, -30, -15, -74, 122, -99, 34, -49, -81, 104, -40, 60, 82, 31, 24, 77, 88, -70, -35, -45, 90, -65, 18, 49, 63, -77, -78, 48, 1, -80, 47, -111, 19, -96, -56, 13, -66, 106, 92, -19, 83, -76, -87, 37, 83, 65, -14, 43, 123, 79, 126, 86, -113, 16, 7, 78, 67, 57, -2, -59, 106, -83, -42, -3, -50, 30, -118, 12, 9, 102, 121, -36, -102, -94, -127, 109, 100, -12, 24, 95, -61, 22, 53, -46, -90, -67, -96, 105, 118, 31, -82, 96, 76, 5, -35, -102, -93, -25, 38, 44, -51, 31, -120, -25, 66, -118, -44, 38, -2, 108, 5, 65, 2, -69, -108, 40, -8, -76, 18, -18, 83, 64, -49, 32, -59, 44, 58, -23, -108, -31, -107, -31, -128, -98, 73, 66, -88, -99, -24, 38, -118, 110, -25, 12, -87, -5, -75, 33, 48, 71, -113, 3, 7, -34, -93, 77, -117, 94, -74, -97, -65, -53, 0, -65, -23, -55, -126, 17, -25, -22, -73, -15, -40, 31, 125, 1, -102, -78, -94, 74, 121, -78, -50, 1, 16, -15, -50, 27, -49, 4, 58, 14, 79, -69, 78, -71, 4, 80, 74, 107, -70, -126, -36, 19, 33, -38, -108, 59, 12, -73, 6, 6, -23, 84, -121, 121, -59, -43, 21, 21, 89, -49, -93, 40, 10, 113, 97, -113, 65, 44, 122, 124, 46, -41, 15, -49, 49, 35, -118, -67, 90, 16, 67, -61, -28, 74, -67, 42, -97, 82, -65, 120, -95, -30, 33, 44, -44, 2, 59, -107, -82, 53, -111, 92, -116, 32, -85, 61, -60, -74, 123, -98, 70, 62, -30, -85, 9, 31, 85, 40, -15, -108, 33, 18, -10, -62, -66, 74, 68, 121, 96, 115, 47, 113, 79, 59, 18, 123, -7, 86, -79, -12, 116, 119, -78, -42, -94, 59, 117, 119, -28, -26, -117, -123, 121, 2, -57, -73, -52, -117, -79, -84, 126, 96, -98, 78, 27, 48, 73, -108, 6, 122, 8, -6, 113, 59, 81, -108, -10, 70, -117, 90, -83, -105, 95, -90, 25, -90, -35, 101, -78, 14, -110, -80, -18, -80, 126, -118, 96, 71, -98, -26, 65, 39, 96, 51, -30, 49, 71, 88, -8, 82, 51, 37, 105, 18, 75, 2, 57, -88, -24, 107, 55, -6, -101, -91, 42, -102, -81, 10, 97, -50, 112, 35, 117, 80, -42, -41, 2, -99, -81, 122, 111, 98, 31, 89, -11, -22, -37, -82, 18, 67, -103, -55, -67, -76, -17, 103, -50, 30, -15, -80, 108, -31, 83, 97, -78, -87, -72, 52, -58, -24, 46, -75, -54, -51, -114, 63, 55, -22, 109, -55, -83, -122, 19, -21, -69, -126, -46, 9, 32, 68, 57, 13, -91, 12, -18, -41, 53, 39, -117, 123, -113, 57, -79, -39, -122, -65, -103, 61, 41, -122, -121, 87, -115, 26, -62, -56, 28, 20, 81, -68, -40, 11, 73, -2, -105, -72, 85, 77, 95, 97, 72, 110, 26, 121, -57, 33, -71, -32, -34, 98, -25, -27, 57, -12, 127, 123, 60, 27, 16, 13, 88, 104, -104, 33, -26, -80, 89, -68, 125, 56, -99, 69, 38, 55, 63, 110, -40, 120, -50, 55, 90, 53, -100, 20, -87, -100, 15, 101, 55, -97, -13, 15, -120, 11, -79, -18, 59, -118, 42, 56, 67, 71, -2, -23, -1, -67, -41, 87, -75, 38, 14, -113, -37, 43, 35, 5, 71, -77, -22, -2, -46, 93, -114, -38, -23, -65, 73, -92, -55, -13, 93, -116, -69, -37, -10, 58, 24, 77, 17, 77, -13, -96, 92, 79, 75, 0, -44, 18, 51, 62, -112, -123, 28, -98, -32, -123, -35, -87, -87, 39, 28, -122, 51, 87, -31, -87, 17, 121, 119, -93, 70, -22, -61, 35, -71, -114, -93, 13, 32, 86, -52, 48, 91, 104, 79, -69, 109, -84, -28, -106, 83, -127, -99, 7, 88, -2, 48, -22, -8, 39, 13, -66, -110, 80, 97, -53, 94, -124, 89, -2, 90, -91, -82, 54, -115, 125, 113, 122, -86, -42, -112, 125, -41, -83, 4, -81, 44, -75, 25, -92, 92, -90, -30, 110, 118, -60, -70, 84, -56, -109, -46, -93, -72, 1, 89, -59, -2, 74, -65, 40, -96, -49, 38, -9, -3, -86, 39, -87, -33, -64, -51, -68, -25, 47, -86, -35, 115, -28, -78, -68, -9, 4, -33, 47, -123, -72, 116, 4, -126, -77, -84, -93, 3, 82, 26, -128, 125, -63, -87, -36, 2, -10, 24, 105, -91, 67, -58, -103, -89, -8, -43, 31, 125, 52, -50, -126, 108, -61, 6, 110, -10, 51, -111, 121, 5, 44, 121, 2, 109, -94, 95, -17, 24, -9, -40, 62, -70, 31, 87, -30, -105, -84, -127, -108, 96, -49, -105, 76, 18, 29, 58, -119, -48, 76, -126, 86, -8, 124, -40, -27, -98, -73, 85, 55, 47, -83, -11, 105, 76, -52, -53, 100, -8, -52, 120, -40, 28, -113, -92, -82, 45, 94, -73, 125, 42, -70, 83, -94, -74, -84, 8, -44, -29, -35, -117, -110, 10, 0, 124, -41, 76, -57, -69, -60, 20, -77, 28, -80, -61, 64, -34, 112, 31, 22, 109, -55, 80, 65, -20, -122, 109, 116, -38, -48, -47, -26, -29, 91, 102, -33, -78, 51, 38, -19, 119, -70, 33, 20, -22, 100, -44, 73, 84, 115, -33, 65, -67, -81, 2, 41, -75, -17, 29, 15, 64, 110, 117, -93, 73, 92, 2, 124, 15, -88, -23, 6, -29, -118, -102, 77, 110, -17, 22, 66, -30, 117, 4, 31, -92, -122, -56, -39, -10, 101, 105, -74, 83, 94, -39, 29, 58, 91, 25, -55, -125, -126, 80, -26, -115, 106, -76, 123, -39, 74, 62, 60, 64, -62, -37, 100, -56, 36, -66, 62, 9, -89, 116, -35, -123, -51, 122, 64, -88, 19, -119, -84, 21, 89, 18, 34, 68, 70, 30, -99, 17, -36, 89, -47, 30, -75, -75, 102, 89, -13, 37, -30, 26, 25, 63, 32, 103, 57, -32, -113, -52, -23, -69, 98, -61, 78, 4, -121, 20, -94, -92, -91, -2, 126, -10, -100, -77, 44, -125, -116, -97, 40, -18, 58, -63, -82, -38, -88, 103, 58, -72, -76, -93, -13, -106, -26, -63, 26, -19, 86, 61, 18, 123, -69, 16, -14, -40, 67, -98, -37, 79, -67, -125, -67, 119, -60, -21, -47, -19, -45, -117, 37, 7, -81, -104, 29, 21, -38, -73, -125, -80, 116, 21, -85, -80, -91, 29, 8, 104, 59, 99, 55, 121, 102, 116, 112, -86, -32, -62, 23, 51, -51, -68, -70, -4, -43, 87, -110, 47, -114, -107, 95, -125, 42, -118, -77, 79, 40, 59, 55, -29, 30, -18, -36, 4, -30, -51, 46, 66, 15, -58, -11, 92, 2, 47, -39, 87, 6, -21, 6, 21, 0, -27, 24, -86, -16, 75, 121, -104, 6, 48, -5, -92, -98, 88, 40, 0, -91, -42, -61, 52, 28, 56, 16, -97, -24, 105, 118, 110, -44, -3, 3, 84, 98, -101, 126, -46, 102, 119, -22, -20, 39, 102, 16, 69, 62, -72, -58, 99, 15, 9, 23, -85, -63, -89, -54, 41, -111, -63, 24, -27, 62, -101, -70, 32, -73, -72, 115, -99, -80, -35, 10, 87, -61, -102, 29, -127, -45, 99, 100, 98, -20, -5, -115, 45, 35, -40, -41, 52, 25, 111, -103, -41, -118, -45, 119, -63, 12, 106, -33, 60, -56, 105, 19, 11, -125, -80, 13, -42, -109, -15, -72, -1, 109, -58, -83, 16, 30, 4, -60, -73, -13, -35, 14, -3, 49, 5, 63, -67, -16, -98, 121, 56, -121, 12, -61, -118, 61, 80, -31, 80, -62, 25, -48, -81, 95, -3, 63, -3, -127, -125, 52, -12, -32, -62, 113, -111, 72, 48, -50, -72, 78, -57, 112, 85, 84, -77, 96, 17, -124, -63, -31, -58, 90, 49, -11, 58, -82, -76, -73, -81, -73, 108, 35, 23, -82, 21, 41, 118, -59, 119, -82, -108, -65, -98, 105, -109, -46, 73, 36, -42, -118, -123, 28, 101, 55, -111, 31, 101, -59, 86, -107, -4, 66, 56, -109, 113, -51, 60, 103, 19, 52, -106, 39, 115, -76, 16, -122, 6, -38, 42, 92, -28, 47, -8, -55, -26, 9, 104, -52, 78, 63, -31, -54, 1, -103, -34, -14, -25, -102, -38, 122, 78, -16, 33, 65, 36, -79, 71, -85, 11, -15, -121, 112, -95, 0, -71, 7, -119, -94, 83, 88, 97, -76, -94, -30, -50, 0, 85, 53, 27, -81, 47, -23, 31, -48, -85, -61, 1, 114, -18, -115, -28, -10, 125, 5, 118, -74, -116, 127, -40, 96, 87, -71, -108, 122, 28, -30, -6, -15, -105, -107, 32, 70, -1, -65, -106, 42, 2, 24, 28, 113, 37, -128, -25, 34, 5, -35, 88, 18, -36, -79, -14, -76, -22, 6, -82, -122, 105, 40, -9, -128, 62, -105, 71, -67, -42, 93, 103, 89, -11, 3, 74, -102, 4, -79, 60, -119, 14, 21, 27, 106, 70, -115, -98, -80, 20, -52, -73, -3, 117, 46, -3, 51, 70, -60, 112, -100, -94, 87, 117, 23, -38, 63, 50, 94, 112, -18, 104, -2, -125, 3, -23, 73, 17, 7, 122, -91, 84, -79, 34, 73, 95, -97, -4, 37, -28, -20, 66, 6, -61, 55, -99, 29, -9, 79, -4, -25, -66, -28, 102, -63, 103, -49, -117, -8, 86, -123, 29, 42, -74, -65, -13, -107, -33, 111, 59, 67, -37, -3, -55, 30, -76, -26, -68, 43, -74, 56, -109, -12, -100, 121, 53, -125, -56, 64, -4, -98, 69, -103, 73, 123, -39, -68, -111, 56, -84, 76, -5, 7, -55, 68, -90, -3, -86, -30, -87, -32, -102, -68, 84, -74, -75, 10, -71, -3, -54, 53, 27, -112, 79, -28, -117, -88, 33, -100, 96, 77, 104, -37, -44, -79, -97, -6, 47, -55, 92, 88, 42, 118, -108, -2, -84, -55, -120, -26, 70, -45, -101, -31, -29, 106, 70, -18, -110, -25, 11, 114, -76, -13, -51, 8, 37, -20, -125, -44, 54, 95, -84, -32, 86, -64, 94, -126, 9, 103, -24, -49, -70, 4, 48, 29, -18, -10, -117, 1, 93, 22, -13, -111, -118, 65, 26, 47, -83, 29, -125, 99, -4, -81, -61, -46, -17, -94, -43, 120, -119, 61, -57, -61, -63, 119, 96, 48, -18, 107, -79, -53, 2, 36, -35, 12, -27, 119, -69, 19, 20, -66, -10, -112, -19, 58, -29, 92, 92, 56, 84, 101, -11, -101, -88, 55, -110, -120, -25, 0, 115, 24, 76, -11, -68, -87, -127, 34, -96, -68, -75, 52, -6, 43, 68, 103, -27, -89, 67, -63, 95, 23, -90, -43, 50, -50, -116, 69, -42, -13, -59, -54, -117, -111, 63, -57, -70, 65, 105, -38, 125, -98, -114, -8, 74, 83, -33, -81, 122, -93, -15, 90, 58, 23, -81, -19, 102, -69, -78, -68, 46, -9, 6, 57, 9, -58, -128, 67, -121, 106, -98, -124, -120, -84, -4, 82, 127, 92, -126, 122, 127, -13, 84, 57, -118, -125, -90, 112, -66, -40, -83, 108, 80, 51, 37, -39, 121, 37, -100, -128, 15, -70, -123, 24, -25, 1, -22, -26, -35, -20, -32, -36, 95, -76, -106, 106, -73, -68, 90, -11, 21, -121, -31, -27, 59, -122, 62, 52, 44, 90, 53, -69, -107, 58, 83, -4, -69, -66, 98, 25, 42, -61, 117, 10, -9, -117, -12, 47, -56, -50, -92, 93, -42, 6, -62, -111, 12, -128, 69, -72, 90, -6, -12, 111, -76, -57, -21, -16, 5, -50, -119, -80, 17, 126, 58, -120, -118, -82, 55, -46, -4, 92, -81, 82, -30, -15, 99, 110, -15, 41, -89, -53, -93, 27, -69, -40, 98, 38, 72, -24, 116, 81, 24, 5, 79, -46, 14, 89, 0, -59, -85, 124, -95, -38, 79, 3, 75, 50, -14, -68, -37, 25, 8, -1, -76, 67, 87, -106, -23, 31, -2, -34, -16, -106, 99, -65, -24, -15, -103, 104, 55, -60, 101, 88, 31, 52, -36, -22, -26, 78, 39, 66, -25, -81, -63, 27, 114, -104, 49, -37, 55, -80, 57, -89, -58, 29, -26, 47, -114, -1, 23, 69, 68, -4, 30, -29, -80, 122, 77, 23, 72, -12, -39, -81, 35, 26, 74, 21, 50, -5, 113, -23, 43, 42, 16, 114, -57, 118, 33, -42, -10, -72, -101, -70, 53, 57, 29, 101, 51, -22, -4, -5, 95, 85, 42, 2, -17, -12, -104, -95, 112, -119, 10, 27, 51, -102, 13, 123, -111, -82, -47, 7, -25, -20, 65, -100, -90, -34, -127, 89, 72, -2, -43, 39, -45, 127, -86, 67, -12, -62, 100, -28, -53, -17, 127, 126, 9, 13, 121, 26, 59, -54, -95, -94, 55, 98, -66, 93, -64, -64, 54, -119, 62, -117, 48, -111, -117, 90, 84, -1, -100, 57, 99, -25, -88, 98, -26, 49, -17, -33, -52, -85, 42, -19, -51, -31, -48, 12, -66, 16, 76, 116, 25, 10, -128, -54, 27, -117, -92, -16, 10, -63, -87, -19, 40, -47, -49, -114, -126, 63, -18, -50, 106, -104, 60, -73, -7, -116, 67, 55, 28, 15, 43, -74, -103, 43, 0, 53, 54, 36, -91, -64, 101, -50, 45, 14, 31, 125, 28, 33, 60, -118, 112, 38, -94, 44, 93, 27, 56, 33, -46, -44, -80, 126, 10, -54, 41, -118, 127, -32, 47, -92, 32, 20, -14, -50, -94, -111, -53, 63, 50, -121, 73, 34, 45, 108, -50, 10, 7, -122, -85, 90, -37, -36, 88, 101, 38, 1, 112, 37, 97, 31, 73, 2, -77, -69, 80, -42, -52, -101, -107, 126, -94, 94, 33, 79, 74, 111, -39, -46, 118, 5, -84, -47, 97, -124, -74, 7, 5, -90, -84, -25, 69, 117, 105, 121, -80, 57, -49, -4, 84, -28, -6, 118, -62, -101, 69, -115, -117, -98, -33, -127, 35, 11, -46, 4, 15, 8, -117, -108, 47, -73, -5, -12, -84, -28, -19, -36, -99, 60, 88, 113, -96, -45, 103, -29, -18, 44, -16, -7, 75, 79, -6, -18, -38, 76, 115, 105, -43, 126, 125, -124, -74, -7, -8, -30, 93, 102, 63, 123, 34, 23, 108, 67, 106, 84, -90, -39, 0, 22, 82, -53, -27, -51, 58, 63, -103, 45, 40, -18, 43, 37, -14, 97, -98, 107, -60, 124, 81, -125, 119, -13, 26, 99, -74, 5, 55, -36, 94, -72, 114, 48, 3, -41, 125, -67, -106, -105, 106, 62, 5, 22, -28, 120, -9, 2, 99, 59, -2, 52, 62, -11, -89, -39, -39, -34, 94, -112, 58, 60, -56, 45, -20, 76, -124, -22, -119, -101, 1, 116, 89, -122, 10, -67, 126, -127, 64, 97, 61, -66, 21, -5, 52, 61, 84, -115, -101, 50, -99, 85, -18, -26, 2, 91, -78, 7, -59, -69, 34, 70, -81, -5, 76, 57, 57, 75, 59, -7, 44, -8, 55, -62, 115, -21, 127, 72, -8, -102, -6, 22, 111, 105, 124, -14, 68, -82, 121, -119, -23, 27, 79, 25, -106, 27, -46, 79, -26, -115, -56, -109, 5, -128, -43, -7, -21, -44, -63, 100, -18, 59, -6, -35, 36, -10, 79, -24, 36, 72, -15, -115, -29, -64, 38, -6, 92, 121, -55, -62, -122, 18, -43, 12, 18, 42, -123, 125, 126, -58, 97, -20, -127, -37, 74, 38, 81, 25, -114, -11, -30, 0, 3, 69, 64, -87, -65, 28, -94, 9, 95, -87, -101, -76, 53, 45, 95, 58, 42, 93, -128, 12, -54, -127, 103, -108, 39, 57, 45, 54, -82, -113, -74, 49, 85, 118, 91, -108, 19, 125, 29, -14, -90, 56, 38, 91, -27, 5, 21, -112, -29, 21, 28, 45, 23, 3, 65, -66, -68, -18, 116, -21, -2, -86, -100, -45, -95, 119, -25, 52, 117, -123, -90, -101, 61, 76, 119, -93, -46, 12, -77, 53, -94, 79, -30, 57, -46, -93, 119, 15, 17, 108, 122, -113, -106, -106, -30, -73, -114, 74, 107, -125, 79, -111, -98, 12, 94, -107, 47, -80, 34, 98, 101, 68, 49, -57, -3, -124, -22, -12, 19, 123, -32, 13, -117, -9, 35, -19, 46, 49, -73, 26, 52, -122, 43, 83, 19, 9, 104, -62, 57, 10, -91, 30, -50, 86, 101, 75, 90, -49, -64, -19, -53, 32, 122, -42, -105, 30, 67, 70, -49, 123, -32, -124, -127, -117, 87, 20, 21, 63, 87, -50, -54, 124, 109, 24, 82, 82, -28, 45, -94, 36, -102, -19, -60, -107, 67, -36, 51, 6, -94, -126, 1, 2, -122, 3, 13, 93, -105, -94, 29, 110, -15, 103, 106, -34, -1, 61, -80, 99, -22, -46, 7, 4, 63, 76, 25, 2, -88, -52, -119, -54, -49, 10, 76, -43, -115, -39, -77, -91, -4, 80, -109, 109, 55, 126, -53, -74, 59, -5, -102, -91, 78, 33, 41, 13, -19, -61, -112, 21, 15, -103, 95, 94, 35, 43, -76, 49, -123, -25, 86, 1, -73, 105, -18, 110, 103, 57, -92, 34, -76, -66, 71, -126, 96, -15, 16, -51, 52, 32, 99, -61, 57, 66, -94, -36, -18, -42, -115, -13, 61, 99, 116, 116, 77, -30, 98, 52, -101, -122, -41, -49, -59, -98, -46, -91, 15, 98, -14, -61, 2, -43, 7, -69, -104, 41, 23, 6, 127, 37, 121, 60, 8, 109, 48, -43, -49, 18, -118, -22, 24, -31, 57, 93, -1, -117, -126, -113, 109, -11, -46, -17, 74, 89, 42, 98, 2, -62, -24, 1, 103, -31, -67, -17, -50, 109, 69, 29, -1, 79, -121, -104, -80, 65, 117, 47, 76, 120, 62, 58, -19, -111, -87, -73, 106, 84, -102, -19, -106, 2, 110, 125, 100, -84, -20, -78, -103, -79, 80, 25, -128, 87, 49, -80, 24, 38, 96, -27, 30, 30, -97, -117, 47, -56, -61, 26, -100, -35, -121, -78, 95, 117, -81, 67, -95, 28, 118, -69, 77, 70, 84, 78, 29, 5, 126, -74, -85, 94, 27, 74, -3, 58, 85, -84, -126, -104, 70, -97, -11, 77, -47, -43, 67, 1, -104, 100, -99, -114, -97, 106, 84, 115, 56, -14, -8, 55, 40, 36, 21, -61, -18, -110, 125, -61, -65, 127, -36, -123, -98, 81, 83, -16, -90, 22, 113, -65, -6, -114, -51, 26, 120, -94, 13, 49, 20, -122, -24, -68, 42, 125, -1, -104, -112, -4, -37, -49, -5, 55, -44, 26, 9, -89, -118, 47, 61, 123, 110, -72, -119, -68, 82, -127, -34, -33, 50, 114, -27, -102, -82, -113, -104, 45, -89, -88, -87, 3, -9, 36, -70, 75, -66, 67, 115, -56, -13, 48, -61, -31, 104, -52, 29, 58, -50, 123, -102, -128, 109, -1, -101, -101, 15, -77, 72, 54, -37, 113, -71, 82, 22, -12, 29, 84, -73, 16, -99, 42, -63, -32, -116, -87, 45, 41, 100, 123, 37, 126, 123, 18, -3, -106, 46, -116, -55, -10, 67, 36, -24, 124, -10, 126, -16, -108, 82, 40, 36, 111, -46, 101, -48, -34, -113, 125, -120, 115, 120, 45, 113, 115, -65, -18, -118, 109, -5, -45, -28, -66, 120, 76, -70, -18, 74, 43, 2, 28, -45, -89, 12, 37, -116, 92, -124, -101, 89, -116, -114, 81, 57, 127, 68, 120, -18, 78, 102, 105, -94, -54, -89, -102, -106, -31, 8, 96, -116, -117, -4, -33, -78, -120, -123, -66, 100, -119, -38, 61, -107, -24, 14, 78, -24, -45, 70, 86, -95, 44, 63, -61, 118, 102, -35, -116, -57, 102, 108, -44, 113, -23, 51, -93, -15, 56, -31, -42, 65, 59, -109, 86, -92, 34, 36, 12, 117, -21, -30, -106, -105, -95, -38, -114, -121, 55, -102, -50, 29, -121, 34, 14, -16, -42, 49, 97, -114, -109, -73, 80, 78, -53, 38, 114, 109, -53, -2, 98, 54, 96, 120, 77, -127, -46, 91, -120, -118, 118, -41, 39, 125, 121, -74, -19, -49, 103, -50, -34, 122, 6, -82, 73, 81, 84, 59, 62, -97, -70, 32, 85, -102, 24, 35, -100, 107, -2, -92, 117, -12, -5, 28, -15, -11, 82, 94, 68, 58, -83, -94, 52, 51, -48, -3, 4, -91, -71, -62, -60, -13, 98, -102, 13, -6, 61, 41, -27, -69, 78, -38, 48, -55, 119, -95, 62, 73, -128, 3, 3, -83, 37, -72, 96, 118, 53, -28, -101, 110, 38, -33, -31, 8, -7, 111, -126, -74, 24, -24, -14, -26, 66, -94, 48, 57, -61, -18, 3, -61, 113, -122, -16, 23, -66, -48, 13, 116, 52, 40, 98, -38, -121, -60, 98, 1, -77, 101, 55, 75, -51, -87, -78, -113, -53, 98, 73, 15, -48, -52, 82, -62, -46, -61, 89, 17, 19, -26, 5, -56, -114, -25, 34, -107, 43, 5, 22, 94, -22, -50, 42, 55, -9, 92, 70, 67, 62, 15, -46, -114, 91, -92, -48, -82, -25, -87, 63, 123, 15, -60, -61, 29, 43, 101, 51, -41, -22, -55, -75, 84, 23, 95, 11, -113, 59, -46, 82, -7, 97, -92, 8, 61, -56, 88, 107, 48, -126, 42, 43, 17, 110, 110, -81, 25, 83, 98, 112, -66, -85, -90, -110, 67, -123, 30, 82, 65, 112, 36, -70, 81, 72, 66, 14, -112, 27, -7, 64, 29, -93, -21, -82, -111, -39, -35, 43, -83, -65, 27, -21, -21, 65, -3, -82, 71, -101, -128, 8, -117, 36, 66, 93, -20, 5, -21, -4, -96, 101, -67, 61, -120, 40, 107, -102, -126, -55, 69, -81, 8, -32, 26, 115, -94, -105, -95, 105, -77, -95, -15, -66, 69, -77, -101, -79, 56, 7, 46, 88, -20, 107, 21, -12, 19, 1, 14, 21, 74, -45, 68, -46, 52, -34, -58, 86, -10, -25, 63, 41, 9, -80, 103, -50, -29, -125, 0, -100, 10, -82, 116, 118, -103, 10, -22, 44, -117, 121, -62, 85, -52, -122, -89, -128, -27, -19, 86, 91, 85, 21, 4, -34, 69, -21, 44, -87, -18, -84, -59, 120, -38, -71, 110, -13, 67, -39, -96, 78, -46, -30, 35, 30, -24, 75, 31, 77, -72, -11, 40, -115, -117, -84, -21, 80, 24, -104, 121, -122, -60, -66, 127, 31, -8, 109, -110, -69, -58, -78, -118, 24, 20, 45, -73, 125, -8, 86, 74, 49, -53, -13, 62, -42, 31, -86, -89, -73, -62, -96, -66, 6, -33, -67, -91, 87, -86, -72, -110, -15, -22, -100, -119, 127, 74, -64, 124, -62, -106, 70, 115, -30, -71, 50, 56, 89, 92, 95, -112, -98, -128, -50, 36, -33, 11, 74, -74, 54, -126, -56, -89, -20, -27, -80, -21, -81, -15, -25, -15, 7, -82, -27, 105, -25, -105, 34, -64, 115, 1, -47, -111, 1, 31, 53, 96, -85, -1, -106, 97, 1, -33, -120, 110, 68, -72, -39, 115, 41, 65, -28, -79, 111, 73, -102, -42, 96, 60, 23, 83, -66, 104, 100, 63, 7, 26, 32, 50, -103, 54, 19, 27, -107, 27, 9, 89, 84, 98, 76, -3, 35, -79, 46, 18, 122, 73, 105, 91, 5, 0, 46, 67, -24, 19, 3, 111, -83, -93, 34, -58, 89, -75, 97, 111, 81, -22, 72, 37, -51, 21, -94, 112, 70, 81, 3, 64, 26, -20, 27, -97, 108, -54, 99, -44, 93, -26, -61, -118, 9, 101, -48, -30, -101, -78, -47, 108, 28, -102, 17, 105, 47, 51, 90, -11, 4, -35, -75, -98, 73, 81, -66, 53, -101, -95, -119, 120, 7, -52, -126, -112, -78, -46, -14, -51, 4, 68, -71, -95, 94, 74, -118, 13, -3, 100, -126, -126, -63, -73, -96, -118, -120, -34, 63, -93, -1, 72, -101, -122, -107, -99, -106, -57, -16, 9, 20, 116, -51, 77, -107, -85, 23, -96, 56, -108, -124, 58, -106, -58, 113, -73, -48, 122, 21, -112, -99, -107, 88, -71, -101, 109, -42, -78, -76, 70, 59, 72, 59, -120, 21, 80, -77, -84, 112, 107, -63, 117, 37, -41, -69, 22, 14, 11, 16, -92, 27, 46, -71, -12, 103, -44, -31, -67, 6, 22, -124, -63, -34, 63, -55, 116, 15, -4, -96, 0, -25, -31, -11, -116, 57, 48, 35, -57, -69, -77, -21, 87, 97, 36, -53, 72, 121, 44, -122, -1, -62, -118, 65, 33, 73, -118, 21, -40, 7, 53, 88, 110, -105, -51, 123, 80, 125, 30, -105, -71, 81, 3, -112, 51, -89, -37, -5, -96, -121, 1, 32, -54, 11, -31, 107, -44, -21, 0, 45, 114, -75, 5, 97, -52, 83, 92, -100, 80, -6, -76, -119, -53, 55, -103, 126, 94, -12, -6, 127, -4, 123, 31, 70, 7, -128, 49, 91, -21, -79, 8, -34, -26, -114, -65, 51, 97, -101, 79, 49, 21, -125, 59, 96, 58, 84, 95, 25, -55, -39, 24, 69, -44, -73, 11, 91, -73, -68, 55, 34, -19, -65, -128, 83, -51, -65, 6, -82, -38, -42, 96, 111, -39, 27, 80, -108, -17, 47, 45, 56, -120, -59, -3, -36, -4, -120, -72, 51, -60, 111, -43, 49, -82, -42, 5, -4, 21, -117, 42, 112, -31, 10, 95, 59, -91, 47, 79, 21, -34, -4, -51, -26, 65, 75, 67, -67, 83, 123, 112, -104, 106, -59, 73, -104, 27, -50, 20, -79, -38, -65, -95, 59, 73, -128, -10, 111, 48, -59, 4, -114, 65, 81, -11, 2, 28, -72, 63, -16, -77, 47, 8, -99, 117, -47, -75, 16, 32, 74, 65, 122, -119, 98, 53, 82, 99, -84, 65, 19, -15, -59, 33, -77, -105, -106, 53, 51, -50, -11, -93, 1, -92, 43, 30, -103, 125, 84, 42, 29, 30, -21, 23, 39, -50, -52, -7, -79, -8, -69, 68, 106, 0, -27, -99, 23, -4, 82, -53, 74, -57, -18, -52, -20, -102, 106, 5, -105, 62, -81, 52, -36, 27, -53, -125, 105, 23, -3, -102, -112, 56, 94, 122, -72, -61, -105, 80, 63, 105, -101, 10, -79, 9, 86, 29, 35, 64, -94, 58, -1, -46, -18, 91, 109, 57, 95, 86, -47, -36, 112, -31, -108, 78, -37, -52, -111, -14, -100, 81, -37, -73, -37, 12, 65, -79, -87, -28, 113, -52, -97, -16, 30, 13, -52, 11, -57, -85, -31, 24, 7, -47, 121, 27, -97, -44, 103, -80, 70, -124, -127, -95, -69, -36, 46, 124, 13, 87, -31, -1, -93, 0, 111, 65, -115, -69, -52, -44, -26, 45, 108, 109, 126, 101, 8, -99, -71, -16, -50, 127, -12, -49, -95, 47, 44, 79, 44, -71, 38, -115, 56, 74, 13, 40, 11, 26, 99, 88, 111, -54, 5, 91, -73, 4, 65, 64, 33, 122, -80, 111, 122, 36, -65, -101, -45, 107, 106, 127, -92, 16, -116, 93, -38, 25, 5, 102, -76, -24, 62, -93, 50, -61, 126, 106, 71, 63, 42, -23, 58, 90, -40, 52, -2, 23, 79, 81, 2, 57, 81, 39, -55, 93, 4, 36, -9, -119, 10, 43, -15, -56, 78, -92, 11, 76, -114, -45, 12, 56, 60, -58, 18, -108, 122, -112, 44, 73, 97, -82, 2, 50, 85, 75, 16, -39, -17, -121, -30, 121, 50, 84, -63, 0, 120, 77, -52, -122, -96, 88, 62, 92, -98, -48, 112, -104, -32, 28, 97, -63, 75, -29, 116, 32, -81, 4, 122, 30, 11, -36, 24, -67, -80, 89, 61, -88, 38, -119, -82, 70, 98, 108, 34, -128, -68, 19, -103, 28, -81, 122, 94, 122, -34, 82, 27, 13, -42, 21, -85, 97, 113, 67, -98, -94, 29, 91, -54, -61, 100, -7, -118, 70, -27, 44, 71, 34, -65, 96, -66, -17, 90, -100, -23, -72, 110, -124, 69, -60, 25, 113, -91, 11, 52, -61, 45, -47, -98, 119, 21, -125, -16, 31, 73, 86, -53, 16, -8, 11, -16, 54, 122, -53, 83, -29, 3, 65, -24, -55, -122, -127, -70, -85, 12, 110, -17, -71, -64, 13, -79, 85, 16, 33, -12, -38, -9, 63, 106, 111, -54, -37, 38, -60, 38, -7, 40, -87, -70, -112, -14, -64, -111, 44, -20, 30, 27, 91, 87, 91, -24, -120, 48, 121, 42, -92, -45, -95, 99, -67, -111, -82, 24, 55, -14, -66, -80, -102, -24, -22, -86, 90, 43, -68, 7, -105, 90, -94, 114, 49, 125, -38, 58, 45, -45, -28, 81, 38, 5, 52, 100, 22, 98, -4, -51, -43, 59, -3, -17, -93, 104, 26, 125, 19, 86, 4, 42, 48, 38, 28, -31, 35, 118, -101, -48, -54, -1, -95, 112, -123, 86, 84, 27, 56, -47, 105, -115, -116, -26, -3, -81, -50, -105, -84, 97, 109, 49, 11, 29, -41, -89, 126, 123, -98, -102, -53, -24, 25, -19, -40, 30, -61, -83, -70, 123, -2, -93, -119, 10, 9, 6, 57, 88, 29, 101, 57, 10, 22, -59, -89, 110, -20, -91, 105, 10, -65, -76, 114, 89, 33, -53, -9, 100, -8, 49, 96, 118, 84, 105, 0, -34, -17, -71, -74, -116, -98, 111, 22, 53, -76, 61, 35, 33, 98, 12, -85, -94, 64, -98, 123, -30, -23, -14, -58, 97, -92, -90, 87, 120, -113, -41, -42, -2, 16, 12, 10, 46, -4, -96, -29, 48, 93, -122, -47, 64, 18, -3, 98, -45, 27, 93, 53, -124, -49, 123, 101, -13, -94, 60, -20, -79, -109, 66, 48, 35, -49, -70, -47, 75, -37, 53, -5, -72, 59, 77, 120, -50, -54, 90, 33, 101, 55, -42, 105, -121, -47, 78, -6, -13, 10, 102, 37, 29, 41, -43, -64, 120, 15, 17, 67, 106, -58, -66, -93, -126, -117, -101, -48, -43, 118, 113, -70, 45, -57, -93, 52, 24, 113, -81, -116, -5, -107, 49, -104, 62, -122, -40, 54, 21, 106, -7, 0, -80, 56, 35, -78, 67, 62, 2, -103, 52, -13, -45, -30, 58, -9, -106, -45, -24, -59, -33, 100, -37, -112, 124, -103, -106, -43, 80, 43, -65, -55, -85, -17, -127, 78, 34, 69, 13, -92, 94, -63, 24, -79, 35, -46, 40, 58, 37, -111, 127, -124, 117, -38, -108, 113, -12, -86, -58, -60, 86, 5, 13, -127, 117, 15, 80, 23, -44, -35, 59, -78, 30, -45, -29, -62, 38, -116, 124, -53, -99, 123, -48, -110, -42, -28, -125, 74, 15, -54, -114, -27, 79, 27, -26, 68, -86, -74, -37, -2, 19, -105, 48, -78, -22, -108, -12, -112, -96, -16, -36, -67, -21, 44, -49, 65, -112, -46, 11, 31, 28, 25, -124, -20, -75, -21, -80, -33, 33, 12, 94, -75, 35, 14, -25, -115, 34, 91, -98, 66, -53, -6, 127, 54, -90, -50, -8, -74, 33, -125, 86, -67, 29, 90, 41, 82, -59, 90, -79, 103, -26, -113, -100, -119, 30, 3, -106, -64, -34, -76, -125, 41, 46, -126, -33, 84, -47, 87, -117, 114, 91, 97, -81, -8, 59, 89, -54, -127, 51, -5, 104, -103, 11, -124, -94, -87, 7, -72, -23, 101, -19, -20, 14, -101, -17, 109, 112, 64, 69, 123, 50, 32, 92, 97, -104, 23, 58, -30, 24, -19, 93, 0, 6, -24, 4, 40, 17, -117, 97, 123, 112, -50, -25, -2, -23, 86, -20, -39, 22, -79, -44, -56, 81, -80, -86, 105, 72, 100, -53, -32, -46, -88, 97, 88, 17, -27, 1, -94, -15, -30, -99, -31, 48, 5, 96, -103, -37, -52, -13, 114, -3, 71, -70, -50, 120, -28, -73, 64, -55, 2, -96, 27, 42, -127, -13, -69, -25, 116, -34, 88, -42, -5, -71, -122, -128, -103, -96, -36, -27, 19, -50, 98, -38, 8, -80, -46, 109, -25, -110, -74, 105, -77, 81, 20, -76, -60, 79, 27, -71, -83, -13, 15, 41, 45, 22, 41, 70, 54, -123, -84, -55, -45, -114, 35, 92, -65, 118, 73, 38, -120, 127, 16, -69, 80, -92, -16, -108, 115, -117, -51, -95, -1, 93, 74, -84, -13, -13, 114, -87, -7, -98, -14, 76, -83, -107, 40, -20, -117, -15, -110, -108, -16, 34, -49, -64, 70, 63, -43, 58, 75, 34, 91, -54, -1, 37, -10, 114, -104, -24, -101, 17, 7, 13, -34, 52, 35, -122, -96, 46, -8, -78, 66, 104, 85, -110, -87, 27, 81, -2, -43, 28, -96, -80, 102, 32, 85, -36, 18, 110, 69, 46, -1, -52, -69, 93, -128, 94, 100, -96, 13, -36, -46, -49, -60, -89, -31, -19, 67, -77, 107, -104, 79, -116, -55, 54, 44, -98, -110, -66, -116, 87, 108, 12, -93, -88, -23, -93, -122, -51, -61, 19, 41, 22, 99, 110, 61, -60, -37, 0, -9, -57, 25, -57, -45, 98, 125, 127, -128, -113, -67, -115, 103, -86, 25, -118, -46, -126, -82, -40, -48, -15, 108, 121, -121, 79, 103, 69, -109, -61, -59, 11, 10, 94, 82, 93, 64, 79, 92, 65, 94, -103, 78, 69, -61, -25, 80, 21, -23, 126, 110, 57, -17, 90, 51, -9, 41, 26, -68, 60, 93, 1, -57, -25, -32, -103, -60, -96, 104, -96, 97, 71, -70, 47, 12, -3, -106, -36, -109, 0, -38, -127, -71, 74, 91, 108, -63, 4, 7, -3, -64, -28, 126, 8, 76, -34, 33, -112, -1, 10, -79, -32, -47, -21, -112, 93, 104, -90, -70, 123, 38, 20, 124, 96, -34, 87, 76, 31, -37, -45, -100, 28, 56, -101, -92, 4, -7, 69, 20, 120, -49, 69, -39, 32, -80, -23, -2, -103, 15, 56, -108, -74, -52, -111, -106, 43, 104, 98, -54, -60, -74, -25, 96, 110, 2, -124, -14, 123, 73, -122, 116, -103, 76, -51, 57, 124, 54, -73, -107, -59, 111, -86, -5, -68, -69, 17, 103, -93, -12, -79, -25, 42, 24, -57, 24, -102, -53, -118, -106, -107, -112, -118, -82, 92, -41, 103, 89, -115, -97, 110, -46, -114, -104, 78, -54, -45, -33, -79, -9, 83, -29, 94, -3, 123, -90, -107, -106, -15, -97, -84, 6, -80, -74, 52, -116, 13, 28, 101, 26, 59, 84, 108, 73, 108, 58, -108, -64, -102, -59, 55, 109, 40, 21, -21, 36, 59, 0, 58, -83, 32, 102, 51, 80, -100, -24, 92, 41, -124, 66, -61, 63, 22, -81, 8, 2, 106, 28, 66, -124, 98, -7, 113, 10, -113, -36, -82, 74, 93, 104, 119, -3, 78, 43, -51, 106, -109, -87, 19, -105, 107, 86, 86, 1, -122, -34, -124, 112, 123, 70, 116, 93, -64, 101, -25, -49, -62, 22, -103, -97, -2, -111, 28, -51, 60, 105, -73, 79, -110, 75, 102, 126, 33, 60, -1, 39, -102, 3, 23, -107, -54, 11, 114, 10, -15, -38, 89, 51, 112, 114, 82, -18, -125, -18, 59, 63, -41, 115, 14, -23, 62, -12, -25, -33, -80, 103, -121, -53, -22, 30, -32, 52, -86, -45, -66, 27, 45, -105, -50, 29, -118, -96, -117, -115, 14, 71, 77, 101, 58, -37, -50, -8, 80, 54, 87, -128, 29, 94, -53, -121, -3, 44, 60, 39, 127, 122, -62, 44, -110, 16, -55, -100, 48, -44, -87, -66, -101, 118, -93, 85, -46, -15, -51, -94, -89, -91, -94, 68, -125, -18, 76, 0, -102, 8, -89, -103, 2, -23, 69, 20, 121, -114, 48, 41, -30, 90, 103, -2, 80, -118, -45, -94, -4, 33, -60, 35, 70, -25, -24, 73, 85, -76, -54, 111, 60, -15, -120, -66, 91, 77, 83, 84, 91, 3, -2, -67, -35, -27, 59, -82, -16, -113, -48, 108, 48, 21, 15, -10, 124, 119, -65, 81, -85, 9, 64, 103, 123, 72, -90, 86, 21, 121, 42, -16, -4, -88, 45, 90, 14, -23, -120, 126, -8, -40, 106, -88, 109, -7, 30, 105, -15, 93, 58, 28, -25, -6, 4, -30, -62, 42, -72, 87, 35, 98, -57, -97, -117, 117, 121, 25, -34, -127, 23, 86, -38, 1, 126, -57, 122, 28, -79, -21, -7, 107, -120, 96, -26, 12, -62, 40, -74, -6, 0, 89, -35, 71, 120, -24, 60, 114, -127, -102, 115, 24, 112, -51, -103, 110, 21, -109, 10, 70, -1, -124, 49, 7, 100, -105, -109, -89, 64, -55, 33, -64, -94, 126, -121, -102, -26, 68, -116, -25, 94, -128, 127, 79, -51, -104, 61, 98, -84, -56, 40, 43, -52, -38, -78, -80, -15, -59, -41, -79, 14, 121, -15, 48, 119, -7, 74, -34, -67, 87, 69, -101, 87, 69, 106, -92, 93, 40, -121, -119, 112, 47, 52, -68, -119, 102, -20, -5, -85, 68, 44, 57, 61, -98, -23, 52, 23, -76, -110, 84, -117, 88, 111, 98, 29, 90, -122, -6, 2, -115, 4, -14, 61, -72, 46, 70, -97, -102, -63, -54, 94, 110, -124, 27, -116, -19, -48, 35, 33, -30, -9, 44, -70, -26, 14, 87, -64, 21, -46, 66, 34, 86, -76, -33, -114, 98, -90, -83, 125, -25, -8, 91, -43, -4, -9, -31, 105, 71, -124, 11, -87, -5, -73, -28, 98, 70, -69, -94, -37, 13, 101, 125, -29, -103, -35, -14, 124, 3, 31, 121, 106, -105, 84, -64, 19, -53, 33, -3, -110, 38, -120, -68, -95, -65, 32, -125, -123, 91, -90, -32, -23, -117, -34, 76, -92, 59, -66, -96, -66, 94, -103, -88, 117, 110, -24, 9, -71, -118, -122, -52, 48, -114, 8, 81, -51, -88, 85, -45, -125, 123, 51, -20, -122, -111, -71, -86, 76, -9, -53, -118, -43, -28, -77, -53, -46, 27, 84, 12, 37, 90, 88, -43, 104, -32, -89, -75, 8, 124, 8, 11, 119, -68, 120, 125, -51, -79, -89, -102, 40, -14, -92, 126, 87, -41, -55, -87, 115, -99, 53, 24, 119, 13, 110, 95, 109, -107, -108, -11, -111, 29, -127, -120, 89, 121, -123, -90, -86, -84, -64, 82, 31, -27, 80, -10, 60, -103, 31, 47, -74, -43, -56, -83, 98, -74, -116, 80, -53, -95, -59, -36, 62, -58, -28, 23, -65, -23, 61, -23, 21, 126, -68, -76, -29, -116, 42, -97, -90, -54, 79, -36, 31, -105, 10, 1, -51, 22, -47, 24, 55, 23, 116, -11, 93, -40, -116, -99, 65, 74, 6, -42, 72, 66, 11, -85, 79, -75, -54, 117, -1, -103, -47, -98, -80, 91, 32, -3, -14, 113, -107, -87, 8, -119, 31, -26, -31, 43, 3, -94, -11, -119, -7, -67, 76, -124, -24, 27, -71, 51, 16, 57, 76, 97, 87, 125, 61, -9, -6, -81, -23, 16, -40, 113, 25, 119, -41, 123, 35, 90, -99, -104, 100, 22, -42, 48, 26, 62, -53, 84, -15, 91, 13, -66, 60, -28, -69, -7, 92, 53, 40, -59, -59, -127, -74, 95, 120, 14, 90, 27, -24, 119, 52, -52, 14, -118, 124, -88, 72, -57, 124, -70, -94, 9, -8, 95, 110, 51, -40, 74, -24, -127, -113, 46, -126, -59, 13, 122, 83, -25, 22, -68, -34, -54, 8, 108, -44, 5, -107, -100, 76, -111, -42, 111, 27, 78, 78, 9, 1, -90, -45, 106, -89, -30, 24, -87, 39, -91, -92, -5, 12, 58, 55, 106, -124, -65, 87, -40, 68, 108, -12, 17, 125, 75, 0, 24, 25, -50, -95, -101, -12, -12, -123, 28, 86, 29, 69, -2, 66, 105, 121, -50, 35, 48, -72, 39, 111, -113, 127, 52, 123, -12, -59, 121, -65, 69, 17, 88, -109, 51, 115, 7, -89, 120, -93, 126, 21, 105, -4, -41, 82, -11, 37, -10, -91, 94, -99, -108, 109, -99, 72, 105, 17, -115, 98, 80, 82, -13, 40, 101, -90, 28, -19, -50, 20, 16, -52, -86, -7, 72, 1, -52, -67, -89, 66, -30, -123, 95, -10, 114, 124, -65, 91, 13, -52, 61, -35, -97, -79, -122, -124, -41, 34, -15, 37, -74, -126, 113, -32, -5, 57, 98, 71, 118, -119, 9, -40, -114, -23, 79, -128, -27, -114, 92, 115, -38, 25, -48, -7, 74, -42, -2, -94, 120, 111, 71, -81, 113, 57, 15, -19, -14, -15, -76, -23, -6, 62, 65, 8, -89, 16, 9, 12, 30, -27, -1, 121, 126, 80, -14, 73, -90, 112, 107, -97, 96, 50, -50, 81, -21, 93, -66, 94, -49, -13, -57, 73, -79, -120, -46, -40, 25, 91, 100, -73, -64, -28, -80, -66, -76, 35, -121, -38, 19, 114, -7, -13, 37, 71, -59, -112, 37, 3, 110, 116, 118, -75, 61, -89, -66, -113, -1, 87, 106, -28, -114, -86, 72, -65, -23, 124, 98, -16, -42, -11, -29, 80, 105, -120, 23, -82, -104, -68, 49, -121, -80, 40, -68, 110, 79, -6, 125, -49, -47, 104, 51, -32, -110, -5, 31, -5, -9, 1, 108, 77, 118, -49, 29, 95, -41, -75, -115, -17, -15, 63, -10, 34, -25, 51, 16, -74, -83, 13, 5, -1, -11, -72, 95, 8, 51, -2, -125, -86, 127, 111, 120, 117, -66, 21, 85, 21, 74, 98, -123, -68, 33, -5, 94, -120, -82, -18, -65, -36, 123, 68, 91, -15, 125, 58, 121, 48, -72, 124, 91, -73, 108, 83, -84, -86, -24, -127, 64, -77, 100, 69, -17, 5, -64, -51, 14, -17, 59, 77, 75, 54, 17, 38, -89, 14, -32, -96, -65, 24, -99, -102, 79, -119, 109, 123, -77, -43, 125, 115, 8, 97, 56, 119, -26, 121, -60, 116, -24, 127, 65, -77, 54, -45, 89, 93, 97, -71, 126, -96, 81, -101, -70, 32, -92, -89, 27, -41, -3, 24, -53, -123, -7, -125, 125, 96, 124, -63, 84, -28, -63, 22, 23, 119, 105, -16, 84, 74, 41, 82, 107, -6, 109, -91, -102, -111, -51, 54, -23, 74, -50, 52, 79, 72, 55, 76, 40, 52, -114, -4, -104, -49, -110, 48, -58, 123, -96, -102, 70, 74, 109, 49, -60, 90, 86, -33, 108, -93, -107, -43, 109, -29, -119, 61, -85, 64, 9, 83, -12, 23, -48, 13, 102, -30, -67, -84, -34, -35, -57, -92, -89, -76, 85, -20, -114, 43, 75, 122, 79, 96, -49, 60, -61, -40, -7, -17, -103, -125, -62, 13, 26, 18, -102, 1, 117, -41, 45, -45, 53, 116, -9, 92, -88, -52, -56, -73, 119, -109, -79, 70, 115, 1, 3, -73, 89, 124, 38, 114, 127, 104, 0, 26, -5, 26, -101, -16, 114, 72, 67, 39, 61, -70, 3, 101, 6, 76, -100, -3, 95, -50, -60, 83, 79, 71, -118, 40, 67, 48, 27, 67, 24, -101, -35, -109, 53, -8, 3, 39, -64, -58, -50, 125, 0, 82, 99, -122, 30, 127, 4, -3, -51, 72, -48, -100, 15, -38, 69, -46, -118, -32, -107, 35, -5, -14, 54, -80, 106, -70, 88, -85, 0, -90, -88, -127, 120, -117, -121, 22, -117, 11, -108, -40, -45, -28, -11, 98, 63, -70, -75, 73, 26, -54, -20, -107, 61, -93, -59, 39, -35, -99, 82, 93, -60, 123, 94, -68, -122, 102, 83, -111, -15, 103, -22, 69, -53, 95, 39, -118, -103, 92, 84, 51, -89, -64, 72, 100, -29, -115, 11, 64, -85, -34, 30, -17, -39, -4, 43, -33, -30, -2, -15, 84, -27, 91, 25, 49, 58, -64, 59, 83, -99, 15, 6, -60, 80, -50, -88, -77, -37, 51, 116, 6, -111, 18, 117, -22, -114, 33, 74, -15, -97, -69, -59, 5, -106, 94, -74, 80, -98, 113, 35, -69, 1, -87, -1, -47, -9, 39, 4, 82, -37, -8, -39, -20, -118, -50, 87, -103, 111, 33, 10, -113, 92, 79, 20, 114, 45, 74, 66, 75, 59, -27, -121, -68, 14, 6, 13, -123, -82, -110, 87, 9, 10, -80, 117, 21, -1, 76, 46, -18, -19, -72, -3, -55, -121, -111, -69, 52, 91, 125, -1, 23, -30, 6, 83, 112, -115, -31, 117, -69, -13, 77, 68, 125, 125, 57, 18, -4, 6, -64, 107, 115, -8, -24, -67, -1, -6, -8, -77, -43, -10, 51, 108, 88, -71, 64, 73, -58, -95, 62, 1, 20, 11, -59, 17, 9, 127, -92, -123, 5, -28, 112, -8, 93, -39, 53, -36, 83, -82, 16, -88, 36, -61, -107, -4, -4, 85, -59, 67, 118, -124, -60, 10, 15, 10, -101, -104, 9, -65, -98, -114, 36, -114, 6, 1, -25, -68, 93, -70, -22, -19, -29, -114, 48, -8, 10, -83, -51, 80, 112, -61, 84, -76, 77, -29, 62, 104, -4, -57, -88, 26, -43, 76, 40, 92, -51, -112, -104, -86, -54, 2, 24, 45, 16, -56, -91, -102, -11, -14, 106, -27, 53, 62, 26, 2, -94, -40, -21, 30, 32, 19, -72, 117, -33, 96, 81, 44, 112, 105, 86, -69, -21, -18, 104, 123, 55, -114, -106, -84, 0, -128, 18, -74, 63, -84, 56, 97, 4, -93, -1, -92, 54, 55, -102, -107, 23, 107, 65, 8, 85, 24, 67, -64, -122, 43, -68, 61, 57, -46, 106, -70, -46, -4, -16, -111, 40, -88, 114, -84, -52, -15, -47, -126, -88, -21, -104, 64, -42, 89, -56, -85, -15, -117, -20, -8, 54, 40, -75, -16, 122, -97, 42, -52, 27, -102, -34, -61, -62, -48, -16, 14, 66, 65, 17, 106, -84, 41, 42, 2, 2, 114, 46, 116, 125, -102, -20, 52, 66, 33, -92, 60, 65, 78, -120, -36, 104, -26, 32, -86, 55, -112, 57, -7, 81, -54, -29, 125, 115, -114, -1, -11, -128, -83, -23, 126, -57, 85, 50, -119, -9, 86, 69, -72, 36, 78, 20, 12, -76, -76, 54, 107, -60, -17, -28, -107, 57, 72, -110, 44, 86, 18, -94, 86, 63, 11, 84, -121, -31, 6, -112, 88, -36, 86, -112, -128, 36, 36, 12, 88, 89, -61, 68, -99, 50, -88, -77, -20, 112, -59, -104, 70, 87, -70, 29, 23, 70, -15, 30, -89, 120, 46, 127, -44, 4, -113, -43, -88, 51, 97, -127, 12, -92, 69, 42, 87, 109, 93, -61, 94, -94, -37, 36, 122, 22, -63, 17, -36, 51, -81, 3, 43, 93, 2, 127, -30, 17, -44, 10, -60, -74, 11, 81, -38, -48, -5, -79, -66, -40, -12, -100, -6, 80, 64, -12, -26, -126, -123, 66, 53, -76, -59, -32, -110, 71, -33, -12, -40, 52, 126, 28, 106, 10, -19, -60, 90, 104, -10, -104, -64, 106, -76, 59, 58, 117, -81, -96, 119, -75, 98, 44, -23, -89, -116, -5, 110, -21, 111, -58, -97, 110, 99, -119, -8, -48, -50, -46, -71, 68, -21, -7, 46, 31, -76, -23, 20, -28, 9, 11, 25, -20, -73, -126, 19, -61, -2, 2, 47, -19, 72, 78, -37, 43, 88, 83, 124, -90, -90, -75, 106, 17, 46, 24, -80, 99, -127, 69, -57, 11, -48, 96, 119, 8, 98, 10, 75, -32, -116, -6, 78, 85, -55, -87, 0, -95, 125, -4, -57, -93, 49, -79, 52, -32, 73, 100, -61, 75, 41, 10, -42, 122, -22, -51, 2, -52, 87, -51, 45, 100, 72, -5, 57, -111, 36, -71, -78, 33, 54, -7, 68, -25, 42, -8, 71, -13, -35, -118, -66, -122, 20, 20, -128, 126, 97, 2, -53, 57, 80, 120, 29, 24, -13, -42, 41, -105, 15, 91, 57, -59, -44, -3, 45, 126, 118, -12, -15, -45, -1, 48, -39, -109, -60, -38, -110, -90, 92, -35, 95, 44, -43, -4, -60, 72, 82, 109, 95, -31, 72, 24, 39, -100, -106, -44, -102, -116, 72, 12, -33, -57, -68, 56, -37, 0, -110, -19, 38, 111, 74, 5, 27, -97, -127, 96, 103, 83, 77, 70, -75, 22, -33, 92, 50, -11, -80, 77, 1, 120, -39, 96, -64, 21, 24, 27, -107, 43, -120, 60, 26, 82, -63, -75, 113, -61, -107, 88, -106, 99, 30, -53, -7, 125, -89, -85, -14, -41, 120, 115, -48, -47, 83, 16, 102, -20, -85, 124, -105, -77, 56, 49, -123, 121, 102, 118, -68, 124, 78, -45, 95, -20, 30, -40, -22, 70, 3, 92, -99, -4, 80, -19, 77, 35, 125, 52, -113, -88, 48, -90, -37, -24, 87, -32, -31, 62, -42, 30, 58, -92, 113, 25, 17, 15, 113, 123, -43, -12, 87, -13, 112, 39, 96, 62, -53, 94, -14, -38, -122, -94, 1, -30, 10, -40, 66, 107, -106, -103, 9, 80, -67, -6, -23, 78, -118, -38, 73, -33, 79, 33, 82, 63, -56, 51, -3, 19, 17, 111, 110, 23, -111, -17, 121, 27, 71, 60, 7, 94, 85, -112, 46, -110, 11, -104, 97, 21, -14, 42, 116, -63, -53, 71, -127, 20, -6, -2, -89, -117, -18, -107, 34, -1, 4, 28, -101, -52, -40, 34, -86, -83, 50, 88, -65, -67, 112, -96, 82, -29, 75, 71, 36, -106, 14, 37, 42, -120, -92, 82, -109, 18, 103, 53, -111, -20, -47, -84, 56, 41, 78, 98, 86, 1, 58, -106, 62, 43, -74, 17, -114, -127, -40, 50, -104, 102, -40, 66, 110, -4, 20, -127, -114, -4, 54, -97, 104, -120, -52, 32, 49, -102, 2, 8, 27, -68, 30, -38, 103, 84, 107, 117, 86, -61, 40, 110, -87, -128, 48, -105, -4, -59, -104, 10, 65, 78, 41, 41, 86, 117, -55, 8, -112, 75, -112, 43, -121, 46, -123, 111, 2, 112, 100, -40, -77, 12, -58, -36, 12, 119, -13, -120, -68, 11, 18, 125, -38, -68, 38, -80, -79, 111, 56, -63, 58, 72, 109, 65, -10, 114, 48, 121, 99, 21, -47, -106, -95, 24, -13, 46, 15, 102, 54, 75, -14, -55, 72, 76, 5, -18, 124, 54, -35, 53, 120, -105, -3, 101, 88, 116, 87, 9, 109, 58, -98, -66, 81, -65, 86, -60, 109, -27, -86, 36, -80, 28, 109, 120, -24, -14, -26, -27, -88, 67, -102, -96, 90, 23, -123, 51, 11, 93, -68, -8, 23, -38, 55, -24, 25, 13, 44, 7, 115, 87, -85, -93, -13, -104, -100, 92, 10, 2, -63, 50, -58, -37, 83, -96, 114, 88, 83, -2, 53, -113, 118, -51, -23, 45, 53, -125, -69, -30, 10, -82, -71, 53, -47, 44, 77, -19, 8, -41, 112, 73, -119, -74, -92, 92, -42, -105, 53, -86, 21, -22, -71, 11, 55, 35, -71, -19, 38, -12, 79, -80, 34, -120, 101, 115, 52, 50, -31, -67, -119, -47, -122, -110, 7, -85, 111, 93, -62, 36, -121, 87, -114, -63, -30, 70, 100, 27, -77, 10, -113, -126, 58, 49, -118, 31, 37, 62, -47, -122, 123, -38, -41, -126, -20, 94, -83, -37, 59, -17, 127, 67, -58, -114, -124, 40, 84, 104, -60, -121, -14, -45, -119, -84, -123, -109, 75, 42, 81, -100, 48, 77, -10, -121, 79, 98, 101, 124, -66, 32, -21, -67, -29, 49, -53, -25, -39, -97, -49, 29, -90, 65, 113, -81, 109, 118, -62, 56, 32, -108, 84, -48, 97, -54, -41, 48, -83, -68, 44, -21, 92, -105, 40, -64, 72, 116, 39, -95, -109, 119, 63, -70, 56, 48, -23, 38, 38, 44, -34, -58, 64, -77, 22, 33, -3, 109, -47, 42, -87, 125, -107, -123, -108, 62, -59, 92, 50, 109, 125, 69, 100, 60, 127, 28, -20, -23, -62, -110, -107, 33, -40, 85, 84, 110, -10, -47, 91, 71, 124, -124, 68, -111, -118, 88, 79, -49, 52, 1, -68, 49, -57, -96, -18, -58, 61, 90, 47, 127, 109, 68, 32, -59, 25, -12, -76, -113, 70, -113, 86, 66, -108, 26, 83, -98, -14, 35, -19, -90, -92, 42, 88, -21, 74, -58, 50, 7, -96, -31, 7, -115, -90, -89, -45, 63, 28, 7, 79, -30, 22, 37, -92, 42, -64, 119, 72, 50, 26, -74, 89, 63, 96, 49, -86, 42, 119, 92, -78, -105, -66, 57, -91, -28, 96, -8, -93, -4, 127, 114, 94, 21, 24, -126, -64, 88, 122, -120, 10, 20, -66, -29, -45, -98, -108, -2, 73, -117, -38, 123, -93, 24, 52, -56, 124, 20, 64, -96, -111, 63, -110, 111, -44, 42, 114, 20, 2, 108, 29, -115, 0, 91, -16, 84, 122, 5, -46, 67, 16, 44, 62, 51, -59, -14, 123, -63, -122, 59, -31, -105, -6, -12, -121, 79, -98, 121, -29, 33, 101, -128, 46, -27, 92, -98, -71, 86, 35, 11, 25, -76, -72, -41, 103, -3, 73, 99, 62, 79, 30, -96, 103, -103, 20, 110, 104, 50, 103, -53, -45, 76, -52, -127, -79, -88, -96, -21, 126, 67, 118, 23, 119, -82, 110, 95, 43, 55, 66, -22, 6, -32, 10, -19, -7, -98, -37, -31, 80, -62, 45, -92, -114, 121, -91, -64, -95, -59, 43, -97, -119, 33, 54, -128, 80, 36, 95, -5, -37, 33, 101, 97, -126, -17, -49, -5, 13, 42, 93, -34, 109, 10, 2, 123, 3, 39, -69, 36, 109, 102, 67, 118, 8, -7, 118, -40, -99, 86, 83, -8, -9, 57, -39, -7, -88, 40, 117, 54, -45, 82, -108, -64, -36, 22, -69, 95, -67, -9, 3, -86, -35, -58, -96, 101, 63, -105, -67, 92, 109, -111, -44, -28, 74, 45, 94, 114, -42, 83, 40, 41, 37, 60, 105, -127, -46, -92, 96, 16, 27, -29, 58, 121, 41, 91, 94, -24, 114, -100, -60, 95, -83, 24, -61, 119, -59, -95, 105, 27, 116, 18, -60, 25, -50, -83, 26, 33, -46, -6, -79, 109, 93, 107, 102, 6, 70, 69, 110, 56, 97, -78, 23, -114, 74, 91, -123, -112, 124, 110, 43, 113, 0, 112, 10, 79, -99, -91, -16, -17, 31, 33, -35, -3, 12, -61, -125, -45, -120, 114, -117, 105, -92, 35, 119, 111, -2, 124, 127, -6, 107, 42, -21, -21, 26, 118, -70, 56, -101, 42, -89, 58, -53, 4, -73, 88, 72, -69, -85, 80, -83, -74, 58, -47, 89, 49, -64, -41, 46, -65, 82, 25, 106, -67, -124, 4, -77, -65, -68, -50, 105, -28, -119, -75, 104, -64, -115, 48, -5, -72, 1, 40, -18, -69, 122, -56, 108, -70, 31, 26, -6, -15, -77, -28, 47, -72, 104, 98, -9, -91, -79, -32, 9, -70, 21, -15, -6, 34, -94, 118, 90, 35, 30, -55, 94, 24, 17, 74, 83, -80, -27, -51, 34, 24, 49, -47, 80, 25, -77, -57, 62, -28, 40, -57, 30, -67, 57, -103, 96, 91, -113, 58, -2, 45, -125, -36, -58, 20, -90, -103, 69, 11, -26, -25, -92, -105, 56, 116, 48, 107, -68, -17, -48, 100, 54, 110, -95, -17, -121, -127, -54, -106, 60, 72, 68, 63, -92, -118, -44, -53, -93, -103, 86, 9, 0, 122, 32, -72, 111, -48, -93, -85, 63, -13, -113, -10, -30, -80, 101, -23, -78, -80, 0, 110, 120, -60, 45, -99, -50, -127, -24, -15, -102, -66, 122, 26, -71, 26, 82, -88, 106, 118, -45, 42, -23, -30, -96, 75, 18, -123, -75, 68, -75, 53, 50, -82, 121, -32, -53, -57, -31, 51, 56, -4, 113, 50, -106, -86, -52, 105, -46, -74, 95, 37, 96, -56, -121, -128, -108, 26, -122, -55, -34, -69, 126, -111, -23, 119, -15, 52, -66, 82, -25, 118, -50, -39, 40, -27, 3, 116, -50, 86, -86, -83, -5, -117, -11, 3, -117, 9, -99, -111, 82, -5, -51, 80, 12, 54, 71, 125, -21, -123, 80, 82, 123, -98, -85, 35, 3, 47, 23, 81, 5, 66, 126, -128, 77, -12, 3, 88, 125, 32, 106, 80, -100, -73, 32, 40, 109, -24, 38, -40, -19, -10, -85, -23, 20, -42, -116, -104, -123, 36, 105, 10, -26, 104, 11, -77, -36, -114, -117, -39, 47, 117, -87, 75, -84, 74, -13, -102, -78, -103, -14, 31, 15, 29, -120, -92, 116, -107, -68, 121, 57, -91, 4, -97, -115, -113, -46, -23, -99, -35, 67, 76, -45, 108, 23, -1, 54, -117, 25, 104, -92, -116, 8, 52, 41, 16, 88, 29, 37, -108, 23, -34, -71, -101, -3, -57, -86, 79, 48, -57, -83, -13, -108, 0, -32, 43, 127, -106, 54, 25, 127, 91, 37, 7, 15, -50, -105, -25, 108, 61, -5, 3, -101, 52, 30, 25, 123, 72, -24, 44, -113, 21, -97, -93, -107, -1, 79, -107, 22, 5, 46, 21, -32, -45, -100, 111, 33, -77, -42, 13, 112, 81, -112, -116, 6, 46, 37, 1, -10, -115, -83, 6, 35, -51, 41, 56, 76, -8, 77, -30, 126, -5, 119, -34, 78, -109, -50, -16, -57, 36, 125, -73, -10, -114, -61, 124, 60, 104, -3, -77, 118, 43, 57, 25, 120, -30, -47, 68, 91, -97, -89, 89, 26, -98, -73, -23, -78, 5, 89, -7, -86, 86, 48, 32, 100, 116, 28, 33, 92, -103, 84, 82, 68, 13, -21, 60, 111, 61, 1, 74, 92, 40, 35, -10, 70, 91, 95, 120, -32, 56, -15, 10, 15, -94, -86, -13, -106, 70, -108, 114, 96, 104, 69, 36, -11, -80, -31, -27, 109, 98, -81, 73, 10, 83, -64, -48, 46, -97, -55, -114, 88, 58, 25, -25, 92, 67, 90, 114, 10, 111, 101, -22, 87, 42, -114, -51, 90, -17, 50, 72, -47, 97, 17, 91, 52, 81, -84, -30, 113, -11, -15, 73, -81, -118, -80, -116, 77, -118, 126, -41, 121, 99, 65, 81, 13, 80, -98, -24, -65, 80, -80, 17, 49, 65, -20, -26, 19, 24, 72, 4, -115, -71, -51, -67, -61, -3, -55, -111, 7, -57, -24, 1, -85, -86, -46, 56, 122, -16, -96, -71, -64, -48, 74, 113, -110, -73, -41, 37, 79, -96, -87, 93, -39, -10, -102, 29, 115, -29, 46, -6, 42, -106, 123, 85, -64, -51, 14, -70, 61, 46, -12, 125, 127, -66, 111, -111, -11, -58, 54, -59, -26, 95, -94, 64, -43, -68, -35, -56, 31, -117, 66, -55, -95, 62, -97, -30, -117, 45, 28, 73, -37, -112, 70, -38, -49, 53, -21, 68, 124, -95, -119, -30, -128, -85, -94, -43, -25, -1, 29, -122, 10, -32, -48, 44, -98, -17, -114, -87, -100, 42, 114, -9, 59, 57, 82, -118, -18, -67, 78, -22, -33, 88, 77, -33, -125, 111, 53, -21, -17, -46, -15, 121, 50, 65, 37, 80, -80, 51, 122, -52, -34, 108, 68, -103, 37, 22, -93, -108, 83, 113, -2, -78, 73, -53, 18, 77, -69, -57, -72, 42, 25, 41, 35, -52, -21, -55, -100, 27, 124, -106, 104, -38, -125, 44, -13, 40, -62, 22, 60, -107, 8, -69, -56, -47, 6, 90, -98, 65, -95, -42, -21, 58, -128, -113, -122, -21, -40, -93, -122, -44, -71, 110, 47, -68, 26, -94, 101, 92, 57, 33, 114, -63, 92, -70, 18, -29, -108, 49, -92, -75, -121, 16, 111, -121, 31, 118, -14, 119, -103, -7, -53, -46, -25, 122, 15, -126, -99, -12, 94, 86, -107, 80, -105, 114, -118, 41, -43, -98, -38, -7, -45, -30, -119, -61, -23, 40, -71, 92, 31, -46, -43, 107, 36, 60, 101, -77, 62, -126, 39, 29, 88, 61, -19, 111, 47, -8, 25, -124, 22, 115, -3, 106, -43, 7, -83, 63, -81, -26, 27, 79, 56, 112, 58, -36, 44, 31, 16, -21, 34, -73, -120, -6, 116, -11, -22, 35, 109, -125, 39, 4, 118, -91, -18, -52, 44, 27, -117, 91, -127, 38, 42, 57, 22, -28, -107, -62, -124, 37, 45, 38, 93, 53, -96, 81, -85, 10, -11, -104, 13, -100, 28, 4, -63, -118, 80, 109, 37, 91, 73, 38, 1, -13, -33, -105, 88, -11, -39, 92, -102, -121, 2, 119, 60, 34, 73, 103, -83, -66, -128, 58, -38, 28, -66, 28, 39, -114, 9, -52, 105, -46, 115, -22, 70, -46, 1, 30, 71, 91, -6, 98, 98, 124, 89, 30, 30, 34, 6, 75, 96, 6, 6, -69, -94, 68, 87, 73, 83, -32, -106, 60, 51, -119, -89, -7, -37, 40, -105, -93, 3, 17, -123, -27, 13, 94, -124, -85, 1, 10, 119, -31, -112, -3, 28, -78, -63, -13, 124, -108, 84, -110, 81, 7, -101, 120, -128, -10, 32, -105, 25, -92, 40, 30, 9, -75, -3, 13, -32, 126, -105, -41, -33, -89, 84, 124, -38, -106, -17, -42, -86, -61, -24, 123, 74, 3, 115, 74, 121, 20, 97, 19, 56, 9, -79, -63, 62, 46, 79, -97, 44, 102, -10, -116, -114, -53, -120, -24, -31, -9, 62, 11, 59, -90, 7, 5, 41, -6, -48, 34, -114, -79, -75, 70, 59, -25, -120, -7, -107, 87, 24, 66, 61, -113, 78, 75, -38, 86, -77, 59, -51, 113, -58, -120, -105, 77, 14, 64, -56, 94, -29, -42, -113, 24, -99, 74, 127, -91, -60, -107, 124, 92, 87, 57, 107, 37, 5, -59, -5, 56, -128, 72, 42, -57, 81, 65, -108, -33, 2, -36, -67, 101, 51, -52, -3, 80, -105, -3, 117, -37, 18, 113, -73, -23, 42, -93, -114, -81, -24, 9, 104, -23, -47, 18, 48, -94, -45, 68, 1, 85, -95, 62, 58, 84, -117, -72, 36, -94, 53, 25, -3, -57, 10, 52, 48, -76, 87, 62, -28, -64, -57, -52, 41, 24, 94, -39, 59, -79, -99, -68, -121, -66, 123, 65, -110, -122, 121, 54, -88, 46, -49, 37, 117, 89, -39, 37, -114, -79, -29, -14, -15, 42, 62, -102, -61, 28, -13, 126, 77, 16, -70, 84, 79, -75, 22, 97, -69, 15, 24, -29, -66, 103, -120, -77, 65, -30, 89, 79, 19, -68, -63, -124, 103, 127, -98, -86, 27, 17, -88, -24, -95, -30, -67, 112, 24, 83, 82, 83, -30, -22, -73, 32, -47, -65, 84, -110, 33, 45, 97, -76, 105, -94, -72, 80, -95, -42, 122, 60, 103, -94, -91, -119, 5, -30, 121, -99, -75, 75, 112, 23, -75, -89, -72, 7, -25, -116, 25, -120, 57, -5, -67, 34, 29, -11, -13, 63, 76, -19, -5, 51, 16, 32, 60, -107, -126, 54, -78, -73, 1, -94, 79, 55, -54, -121, -66, 49, -109, 87, 57, 76, -46, 118, -18, 112, -20, 97, 47, -72, -49, -86, 107, 95, 75, 40, 116, 77, -34, -90, -123, 95, -56, 84, 22, 18, 91, 84, -61, 110, 44, 125, 58, 126, 115, -88, 110, -33, -118, 29, 23, -39, 72, 3, -72, 19, -85, -84, -32, 9, -46, -27, -24, 26, -71, 127, -83, -108, 83, -16, -126, -1, -19, 60, -2, -31, 101, -20, 64, 111, -118, -40, -56, 82, 91, 0, -27, -122, 44, 69, 15, 126, -85, 119, 24, -28, 118, 69, -7, 74, -74, -5, -55, 35, -72, 71, -124, -99, -76, 69, -116, -66, -99, -44, -112, 120, 84, -11, 126, 0, -70, 13, -2, -27, 4, -106, 74, -5, 92, -61, -59, -110, 62, 14, 53, 118, -42, 58, -109, 10, -1, -97, 72, 28, -13, 88, 20, -57, -51, 18, 71, 7, -97, -59, 109, 35, -36, 55, -98, -72, 122, -29, -54, 56, 114, 127, 47, -56, 57, 66, 82, -72, 98, 26, 84, -43, -14, -24, 29, 63, 122, -28, -58, -103, 42, -77, 61, -122, 106, 91, -66, 100, -65, 8, 29, -79, 7, -52, -7, -63, -114, -53, -7, 112, 101, -50, -58, -41, 54, 99, -106, 49, -57, -36, 74, 113, 16, 7, 119, -6, -29, -75, -33, 34, 61, 124, 83, -59, -56, -52, 6, -42, 23, 127, -57, -4, -51, 13, 83, -124, -16, 105, 53, 55, -59, -1, 41, 85, -121, 32, -48, -22, 86, 47, -116, 19, 43, 95, 88, 115, -85, -34, -55, 66, -34, 16, -66, 43, -99, -111, 47, 13, 122, -28, -59, -65, 100, 110, -107, 107, 14, -27, -43, -28, -108, -31, 120, 63, -64, 80, 50, -21, -81, 123, -83, 13, 12, -21, -72, 41, -4, 104, -73, -10, -52, -4, 53, -80, -22, 74, -101, 120, -81, -16, -35, -61, 81, -43, -126, -111, -91, 52, -4, -44, 48, 41, 97, -68, -108, -102, 101, 16, -126, -100, -122, -50, 24, 60, -1, -126, 6, 26, 123, 54, -117, -40, 121, 92, 45, 124, 110, 82, 48, -22, -89, -32, -108, -120, 28, -88, -94, 2, 57, -92, 30, 63, -13, -73, -5, 114, -71, -126, 12, -76, 56, 23, 12, 49, -12, -71, 45, -30, -116, -34, 76, -77, 62, 96, -69, -37, -119, -34, 93, 66, 2, -5, 1, 117, 50, 125, 103, 108, 127, -12, -96, 55, -117, 45, -24, -1, 102, -106, 97, 114, -12, 46, -91, -78, 14, -31, 13, 23, 63, -22, -39, -63, 102, 91, -73, 24, 88, -98, 4, 87, 18, 37, 14, 30, -46, 118, -99, -72, -116, 127, -85, 0, 45, -48, 51, -69, 49, -64, 83, -16, 43, -84, 50, 17, -121, 105, -87, 95, -121, 46, 54, 26, -45, -60, -72, 37, -69, -43, 93, -57, -44, -120, 72, -127, -39, -5, -67, -118, 59, -112, -5, -26, -68, -83, 119, -60, -106, -95, -93, -99, 79, 90, 55, -94, -98, 111, 71, -39, -59, 36, 33, 25, 45, -23, 27, -122, 100, 88, -112, 31, 104, 11, -122, -92, 56, 125, -24, 78, -98, 12, 108, 109, -26, 35, -113, 4, 19, 86, 94, 88, -5, -1, -15, -88, 104, -116, -82, 76, 100, -66, -21, 76, 74, -15, 113, 2, -17, -39, -47, 13, 101, -67, -5, -53, 96, 10, 80, -13, -31, 46, -53, 92, -83, 61, -124, -107, 73, -78, 97, 46, -16, -52, -6, -70, 62, -21, 61, -83, 69, -114, 58, 42, -53, -75, 118, -85, 64, 70, 31, -95, -12, 106, 125, 33, 39, -127, 54, -15, -77, 23, -97, 35, 99, 25, 94, 33, -123, 27, 78, 74, 41, 9, -12, 116, 62, -22, -97, -2, -80, 62, 31, 36, 41, 28, -59, -48, 29, 123, 65, 80, 18, 96, -12, -10, -6, -46, -105, -1, 109, 102, -55, 22, -17, 61, 10, -83, -88, 41, 44, -40, -24, -53, 125, -111, 104, -62, -31, 5, -66, -93, -42, 80, -125, 74, -58, -3, -100, -34, 124, -119, -60, -59, 31, 51, -125, -87, 96, -85, 82, 12, 3, -70, 88, 0, -53, 64, 67, 45, -59, -127, 80, 27, 81, 83, -27, -104, -47, 1, -10, -51, 10, 58, 19, -87, -19, 22, -46, -51, 65, -91, 90, -60, -33, 50, 69, 43, -14, 8, -40, 55, 9, -88, -45, -38, 123, 56, -14, -52, -70, 104, 26, 68, 34, -83, 110, -113, 67, -64, -35, 4, -27, -73, 72, 69, 105, 13, -16, -37, -107, 72, -110, 30, 112, -27, 121, 107, -98, -21, -72, -40, -44, 82, -100, 118, 127, -118, -122, 66, -53, -29, -58, 48, 26, -114, -11, 3, 28, 101, 94, 49, 45, 112, -48, 29, -42, -55, 9, -12, 52, 65, 76, -120, 19, 104, 127, 18, 115, -123, -44, -66, -24, 26, 110, -126, 40, -28, 5, -60, -55, -29, 118, 119, -45, -58, 20, 41, 15, -99, -99, -61, 94, 105, -52, -15, 82, -53, -125, 69, -48, -41, -125, 56, 113, 113, 58, 26, -43, -65, 94, 31, 34, 84, 22, 117, -102, -86, 31, 41, -56, 60, 109, -90, 38, -71, 24, -8, 4, 27, -67, 84, 115, -64, 12, 100, -79, -58, -2, 7, 5, -35, -90, -89, -79, 60, -100, -52, 102, 59, 117, -82, -8, 98, -43, -98, -101, 109, 22, 31, 8, 83, -13, -5, -109, 127, -32, -60, -59, 94, 75, 74, -69, 113, 113, -19, 45, -114, 57, 20, 73, 46, 66, -63, 17, -105, -33, 44, -124, 117, -52, 13, 72, 63, -120, 91, 63, -24, -96, -124, -57, 107, 79, 2, 93, 64, 111, 10, 78, 40, -98, 24, -41, 97, 89, 104, 120, -71, 20, 125, -82, 96, 10, 119, 32, 18, 82, -33, 123, 114, -29, -62, 94, -78, 68, 59, 115, 52, -59, 65, -36, -28, -39, 51, -59, -77, 27, -67, -20, -80, -70, 26, -112, 68, 17, 48, -41, -28, -113, -46, -42, -13, 20, -76, 37, -40, 111, 24, -116, -75, -38, -23, 25, 51, -100, 94, 102, 56, -101, -46, 104, -42, 109, 120, -102, -2, 41, -15, 98, 56, 67, -71, -85, -41, -19, 81, 48, -35, -23, 60, 18, 67, -91, -85, -9, -62, -119, -35, 122, -92, 48, 98, -6, 29, 90, 21, -101, 3, -122, 126, -68, 74, -73, -25, -95, 36, -72, 81, -127, 34, 14, 19, -27, 51, 62, 92, 117, 71, -70, 111, 108, 106, 81, -26, 7, 44, 123, 34, -81, -126, 32, -21, 76, 87, 83, 109, -4, -117, 63, -3, 45, -51, -111, -109, -128, 79, 111, 118, 23, -87, 101, 3, -109, 55, 105, 26, -29, 101, -67, 18, 103, 93, 126, 51, 53, 81, 32, -79, 92, -33, 46, 10, 44, 63, 29, 45, 15, 12, 35, -90, 54, 8, 41, 73, -65, 18, -28, 34, -9, 33, -75, -34, -2, -77, -111, -77, -124, 50, -28, 96, -111, -109, -22, 62, 82, -121, -21, -31, 20, -114, 7, -54, 22, -80, -109, 86, 67, -9, -8, -70, -104, 45, 25, 23, 96, 42, 74, 100, -36, -81, 69, -18, -62, -81, -84, -108, -73, 23, -10, 75, 37, 125, -107, -69, -82, -88, -111, 113, 32, 10, -85, 56, -73, 68, -49, -104, -17, -102, 124, 75, -55, 65, -71, 11, 113, -27, 31, -88, 124, -107, 115, 33, -109, -120, 93, -63, -80, 110, -78, 80, -8, -35, 9, 48, -94, 88, 72, 17, 114, 68, -36, -69, 6, 22, 70, -9, 123, -26, 31, 120, -5, 18, 25, 14, 26, -10, 79, 74, -27, -127, 27, 93, -33, -92, 13, 1, 124, -43, -110, 111, -102, -18, -86, 32, -124, 113, -105, -128, -41, 54, 120, 82, -56, 17, -31, 98, -120, -80, 44, -19, -78, -57, -54, 17, -21, 88, -110, -24, -83, -92, -41, -57, 18, 1, 103, 23, -14, 126, 23, 73, 52, 15, 28, 124, -96, 125, 94, -88, -83, 11, 21, -33, 82, 96, 112, -66, 56, -126, 38, 101, -90, 125, -83, 57, -2, -108, -48, 113, -109, 103, 58, 71, -10, -42, 68, 22, -45, 34, 63, 1, -83, -44, 96, -128, -76, 81, -66, 108, 83, 100, 82, 122, 97, 127, 51, -33, -109, -125, -48, -90, 106, -117, 110, -32, -31, 50, 118, 53, -44, 53, -74, 2, -118, -106, 2, -66, 103, 64, -85, 59, 36, 125, 53, 5, 124, -24, 100, -113, -21, -75, -74, -43, -64, -92, 53, 33, 86, 43, -42, -86, -31, 12, 44, -21, 35, -82, 41, 10, 110, 84, -59, 18, 81, 122, -105, 77, -30, 124, 93, 77, -79, -109, -94, -15, -73, 87, -110, -115, 3, -23, -73, 100, 117, 100, -49, 24, -110, 120, -93, -127, 77, -24, 19, 30, -29, 43, -20, 69, 39, -55, 19, 88, -36, 53, -55, 19, 13, -37, 32, -112, 68, 87, 116, 58, 59, -61, -46, 78, -69, -11, 79, -120, 94, -30, 39, -63, -115, -109, -122, 52, -36, 25, 12, 56, -49, 85, -53, 92, -79, 107, 108, 117, 66, 96, 47, -2, -93, -126, -52, -34, -9, -101, -25, -43, -3, -114, 22, 11, -95, 29, -65, -3, -74, 76, -75, 5, 33, 0, -31, 82, -21, -51, 72, -83, -83, -9, 43, -48, -7, 119, 47, 113, -110, -106, -58, 16, -92, 93, -101, -59, -6, -38, 66, 48, -90, 119, -74, 72, -9, 23, 26, 98, 101, -30, -113, -110, 90, 59, -29, -45, 50, -110, -60, 69, -88, 11, -43, -52, -24, -16, 17, 98, 74, -45, 18, 113, -54, 72, 57, 65, -32, -45, 35, -59, 54, 50, -41, 16, -19, 58, 99, -96, 76, -88, 101, 116, 51, -70, -64, -101, 42, 81, 125, -12, -92, 15, -27, -18, -40, -98, -81, 56, -14, 82, 125, -88, 5, -44, 56, 114, -113, 27, -110, 91, 67, 119, 80, -10, -79, -112, 17, 91, 98, 14, -48, -122, -98, 53, -11, -10, 84, 36, -82, -58, -9, -85, -18, 124, -1, -90, 110, 14, 65, -127, -22, 5, 120, -70, 123, -86, -54, 13, -123, -84, -101, -43, -77, -71, -117, 40, 47, 95, -52, 93, -91, 67, -120, 19, 63, 8, 57, 46, -106, -6, 47, 0, 127, 39, 58, 123, 81, -123, 8, 87, -79, 35, -84, -28, 93, -73, -116, 12, -106, -39, -22, -69, -100, -14, 78, 92, 122, 7, 10, -111, -126, -71, 17, -127, 96, -52, 124, 50, -47, 4, 9, 2, -88, 53, 103, -123, 109, 115, 17, -125, -52, 123, -65, -23, -18, -115, -59, -24, 21, 79, -7, 23, -120, -117, 24, 104, -41, 21, 26, 40, -103, -93, -86, -63, 89, -111, -58, 70, -123, 88, 73, -47, 83, -120, 58, -63, -106, 127, 42, 43, 78, -93, -62, 86, -82, 90, 63, 5, -17, -39, -83, 9, -3, -40, 74, -42, -23, -111, -100, -18, 105, 101, 64, 60, 110, -6, 126, -124, -6, 40, 47, -56, 75, 113, -97, 122, 75, 94, -1, -69, -73, 45, 68, 52, -123, 14, -118, -18, 31, -90, 93, 8, -116, 29, -59, 122, -105, -61, 126, 17, 107, 45, 90, 54, 30, 121, 48, -23, 87, -80, 36, -114, 93, -24, 67, 98, 119, 77, -48, 22, 116, -83, -97, -128, 74, -28, 122, 98, 39, 120, -13, 18, 37, -51, -56, -61, -58, 121, 44, -99, -87, -47, -84, -122, 57, 111, 104, 48, 60, -72, -57, 48, -26, -26, 48, -80, 74, 42, -110, -15, 34, 6, -125, -57, 83, -53, 10, -102, -60, -73, -73, -19, 8, -29, -13, -63, -46, -37, 114, -113, 20, -71, 63, 122, 31, -16, -86, -23, -102, -67, 90, 61, 67, 93, -124, 22, -88, 15, 48, -19, 70, 104, 90, -50, -53, -50, 15, 30, 41, 1, 45, -67, 58, -20, -73, -39, 92, -30, 66, 119, 31, 28, 52, -30, -7, 56, 120, 34, -57, 41, -113, -115, 17, 105, -37, 92, -73, 107, -6, 97, -20, -89, -98, -89, 20, -42, 0, -16, 56, -61, -25, -41, 95, -101, 57, -39, 84, 49, 123, -101, -38, -118, -87, 107, 115, 4, 72, -85, -17, -62, -116, 92, -22, -86, -125, 126, 0, 3, -18, -72, 70, 86, 15, 38, 113, -56, 127, 69, 122, 122, 97, -44, -124, -118, -64, 119, 14, -120, -94, 126, -54, -82, 90, 52, -39, 93, 50, 89, -32, -95, -110, -89, 119, 33, 77, 104, 106, 76, 46, 100, 70, 15, -72, 74, 25, -8, 65, -89, 0, 100, -91, 75, -110, 127, -1, -21, 92, -78, -59, -67, -45, -41, -28, -54, 120, -79, -78, 98, 125, 96, 70, 67, -17, 127, 13, -120, -9, -50, -80, 120, -78, -43, 67, -59, -43, -62, 48, -79, -12, 117, -18, 71, -52, 82, -111, -59, -125, -60, -89, -128, -92, 110, 67, 20, 109, -48, 28, -28, 31, 76, -36, 81, -94, -97, -106, -9, -30, 71, 40, 86, 60, -105, 30, -119, 105, 47, -50, 109, 115, -11, 109, -104, -29, 49, 44, -48, -127, -56, 53, 32, -107, -111, -14, -73, -79, 8, 46, 19, -49, -42, -23, -116, -19, -121, -107, -41, 55, -29, -60, 42, 88, -79, 66, -68, 98, -18, 12, 100, 55, -63, 4, 76, -45, 118, -125, 4, -1, 49, -105, 78, -121, 0, 90, -11, 8, 111, 76, -65, -46, -112, 105, -85, -63, 44, -25, -92, -102, 115, -120, 81, -75, 12, 29, 8, 3, 32, -116, -126, -47, -93, 80, -39, 35, 43, 78, -85, 26, 26, -22, 109, 42, -44, -104, 107, -128, -1, -113, -102, -14, -105, 108, 39, 36, 9, -81, -89, -86, -69, -87, -5, -34, 121, 84, -126, 36, 34, -83, -65, -68, 24, -84, 102, 108, -60, 82, 108, 67, 97, -122, -75, 121, 114, 93, 29, -4, -116, 68, 38, -56, 109, -95, 38, 102, 118, 40, 11, 24, 86, 74, 85, -18, 118, 59, -38, -70, 13, -58, 125, -17, -52, -78, -24, -65, -113, -123, 59, -100, 73, -31, -28, 54, 2, -118, 28, -8, 51, -89, -111, 9, 113, 102, 119, 103, 33, -47, -95, -81, 23, -98, 30, 99, -47, -122, -94, -32, -117, 93, -4, 84, -66, 96, 10, 65, 107, -90, -71, 30, -50, -54, -89, -65, -80, -98, -89, 82, -17, -56, -127, -122, -25, 31, 105, 56, 37, -116, -104, 48, 105, 21, 4, -88, -11, -114, 105, -32, -76, -94, 126, 2, -19, -91, 66, 29, -61, 105, -17, 50, -79, -16, 56, 24, -113, 34, -48, 52, 46, -23, -28, 23, 126, 104, 63, -13, 118, 40, 84, -85, 75, 82, 45, -72, 120, -17, 85, -69, -40, -59, 110, 10, 53, 38, -94, 69, -56, -13, -7, 118, 92, 94, 14, 90, 70, -51, -51, 61, 118, -95, 104, 65, 116, 21, 121, 108, -123, 78, -89, -35, -109, -107, 103, 73, 60, -118, 14, -124, -3, -121, 123, -39, 101, 9, -77, 44, 86, 0, -23, 76, 34, -47, 13, 22, 102, 6, 2, 107, -43, 41, -55, -24, 63, -80, -79, -5, -70, 63, -1, 55, 71, -6, -112, 44, -125, -61, -40, 90, 68, 65, 38, -26, -110, -76, 124, 121, 58, -2, 100, -113, -89, -83, -8, 102, -34, 41, -31, 24, -23, 97, -48, -80, -37, -32, 92, -33, 36, -75, -71, -24, 118, 95, 78, -119, -109, 74, -126, 78, -56, 102, 93, -17, -108, -43, -42, -14, 127, 55, -118, -24, 24, -38, 24, 116, 59, -12, -45, -33, 41, 12, 71, 32, -21, 21, 41, -1, -33, 43, -51, 39, 17, -86, -106, 37, 0, -20, -105, -1, -92, -94, 103, 60, -4, -1, 48, -73, 115, -125, 22, 29, 15, -35, -67, 123, 114, 102, -6, -47, 17, 71, 120, -94, 113, -113, 72, -15, -5, 95, 112, 31, -127, 87, -36, -2, -42, -116, 53, -54, -112, -52, 103, 31, 41, -92, 26, 28, -118, -108, 109, 27, 91, 102, 61, 77, 117, 5, -66, -16, -27, -81, -112, -26, -122, -20, 100, -35, -8, 26, 39, 8, 102, 14, -88, 15, 50, 66, -85, 60, 87, -103, -41, 50, 127, -108, -1, 116, 26, 62, -28, 127, 109, -12, -27, 115, 96, -54, -48, -39, 100, 119, 97, 74, 5, -119, -39, -73, 76, 5, 115, 35, 30, -54, -43, 29, -33, 85, 17, 121, 19, 117, 120, 0, -22, -35, -13, -54, 39, 68, 35, 11, 59, 5, -43, -63, 14, 47, -8, -38, -76, -20, 125, 82, 54, -45, -17, -107, -88, -128, -114, 59, 117, -122, -69, -33, -28, 46, 42, -117, -14, -51, 23, -82, 82, 108, -17, -31, 27, 103, 59, 79, -45, 57, 33, -118, -116, -112, -97, -76, -112, -82, 111, -122, -76, -86, -27, 24, 88, -113, 36, -53, -35, -69, -7, -81, -89, 104, 16, 67, 79, -52, 18, -93, -123, -76, -83, -111, -60, -52, -59, -43, -6, -76, -37, 47, -34, 64, -57, -74, 80, 107, 1, -83, -90, 122, -36, -50, 98, 109, -111, 50, -71, 35, 85, -66, 87, -126, -49, -100, -50, 20, -15, 73, 72, 76, -8, -90, 12, 63, -36, -36, 43, 94, 9, 81, 88, 102, -97, 59, 83, -80, -19, -116, 84, -62, -54, 43, -60, 25, 71, 18, -83, -72, -37, 117, -124, 83, -101, 17, 19, -9, 109, -66, -43, -9, -113, -82, -35, -81, 105, -80, -33, -42, -68, -77, 24, 6, 95, 92, -97, 38, -18, -52, 95, 74, -63, 99, 29, -36, -12, -80, 83, -30, -18, -87, 89, -2, -41, -74, 45, -64, -26, -116, 22, 34, -64, -82, -88, -97, -118, -57, 69, -8, 19, 36, -62, 84, 8, 96, -80, 124, -112, -125, -34, -1, -84, -73, 125, 3, -19, 42, 67, 83, 54, -39, -11, 118, 7, 29, -107, 17, 100, 91, -118, -9, -1, -52, -53, -121, -84, -5, -124, -67, -1, -30, 60, 43, 26, 57, -81, -121, -29, 114, 91, -103, -52, -48, -112, 83, 110, -91, -27, 82, -128, -17, -54, 0, 59, 21, 7, 104, -111, 11, -91, 16, 110, 97, -69, 8, 26, -22, 15, 125, -35, -22, -106, 41, 59, -90, -4, 41, -52, 97, -5, -52, -48, 69, 76, -116, -37, -44, 116, -20, 95, -103, 124, 77, 122, -73, -43, 20, 34, 101, 17, 127, -49, 39, 40, -118, 78, -92, 51, -102, -122, -81, -26, -42, 116, -77, -30, -49, 7, -42, 59, -26, -17, 55, -76, -23, 111, 9, 125, 17, -18, 14, 16, 62, -74, -72, 72, -124, -36, -4, -98, -30, 43, 4, 57, 31, 55, -101, 111, -66, -14, 42, 37, 97, -30, 89, -53, -47, -30, -56, 98, 81, 87, -14, 15, -115, 42, -41, -111, -122, 83, -81, -23, -2, 51, -94, -98, -21, -67, -115, 41, 47, 55, -50, 17, -103, -89, 92, -22, 10, -92, -52, -37, 123, 62, 106, -120, -24, -63, -103, -17, -107, -56, 88, 19, 124, 122, 49, -25, -73, 62, -112, 103, -10, -33, -8, 15, 6, -44, 122, -112, -8, -58, -21, -12, -123, -43, -4, -19, 23, 22, 92, 44, 94, 52, -65, 90, 46, 113, -63, 102, 47, -46, 77, -91, 49, -59, 53, -73, 25, 47, -56, -111, 117, 51, 5, 122, -119, -126, -24, 32, 24, -60, -52, -10, 121, 11, -47, 39, -4, 18, 13, -84, 100, -38, -47, 21, 31, -122, 77, -72, 53, -107, -54, 43, 72, 79, 37, 81, 81, -115, -15, -23, -46, 61, 96, -53, -55, -79, 114, 69, 67, 0, 113, 40, 90, -61, -67, -6, -55, -118, 50, 127, -97, 124, 42, 104, 76, -49, 57, 29, -35, -85, -121, 47, 104, 103, 122, -79, -104, 108, 119, 91, -20, 104, 3, -57, -85, 65, 65, -11, 75, -13, -12, 107, -16, -98, 83, -68, -19, 12, 89, 74, 55, 96, -7, 32, 71, -13, 81, 95, -32, 72, 59, 76, 49, -66, -109, 92, 127, 84, -47, 75, -56, 69, 54, 56, 99, 9, 116, -47, -107, 77, -101, 77, 46, 21, -19, -11, -120, -66, -43, -24, -121, -112, -75, 56, -50, -56, 20, -50, -99, 102, -103, -27, 43, 79, -99, 15, -40, -111, 96, -19, 94, 123, -70, 12, 16, 39, -126, 25, 102, -41, -127, 109, -25, -74, 37, 53, -1, -71, -125, 28, -97, -100, -127, 75, 107, -98, -38, -61, -81, -70, 49, -115, -75, 107, 26, 70, 19, 28, -33, -7, 115, -32, -26, -38, 23, -117, -113, -106, -60, -109, 50, -28, -81, 51, -81, -101, 81, 9, -34, -128, 67, -113, -115, 120, 123, 39, 62, 14, -61, -99, -121, -74, -2, -19, 16, -107, -8, 32, -85, 60, 51, 93, -96, 98, 16, -49, 125, -31, 88, -36, -31, 27, -21, -18, 20, -26, -106, -46, 116, -39, -16, 123, 16, 110, -24, -96, -125, 96, 64, -82, 29, -13, -117, 61, -42, 27, -115, -45, 124, 101, 47, -35, 1, -101, 75, -107, 1, 97, -25, -10, -69, 87, -15, 75, 69, 90, 107, 72, 58, 44, 118, -41, -97, -127, -107, -11, 28, -94, 73, 24, -121, -8, 117, 8, 19, 65, 29, -107, 34, -123, 11, 93, 92, 124, 40, 34, 86, 20, -22, 17, -64, -31, 104, -33, -30, 125, 85, 127, -97, 30, 23, -89, -106, 13, 47, 42, -50, -51, 63, 112, -46, -54, 78, -82, -58, -10, 80, -99, -118, -69, 46, -54, 28, 22, 42, 126, 20, -1, 125, 51, -99, 21, 90, -77, -94, 10, 93, -16, 87, 28, -32, -87, 102, -82, -41, -83, 37, -88, -54, 47, -29, 120, 122, 127, 14, 36, 125, -94, -93, 123, 86, -64, 16, 48, -13, 50, -70, -47, -94, -111, 109, 2, -70, 84, 49, 18, -127, -42, 58, -53, -123, -99, -61, 127, -100, 81, 35, -103, 116, 70, -108, 74, -122, 36, -6, -6, -42, 53, 75, -8, 70, 56, 123, -127, 12, 44, 19, 13, -126, -51, 88, -121, -22, -101, -121, 6, 109, 42, 31, 97, -15, 52, 43, -9, -40, -91, 113, 47, 90, 60, -89, 33, -11, -94, 34, -127, 78, -75, 15, 80, 2, -25, 88, 108, 3, 95, -14, -16, 9, -111, -47, 122, 69, 124, -14, -98, -95, -29, 77, 124, -96, 116, 29, 21, -105, -65, 22, 101, -12, -91, 54, 118, 13, 14, 98, -112, -19, -44, 0, 118, -27, 81, 113, -85, 77, -29, -55, 110, 70, -106, 106, 102, -118, 7, -5, -95, 70, -110, -121, -70, -73, 61, -80, 68, -53, -110, 84, 56, -26, -44, 46, 76, -91, 31, 119, 114, -126, -64, 97, 73, -42, 75, 47, -32, -45, -85, 2, -103, -67, 9, -44, -12, -58, 4, -71, 17, 23, -115, -55, 125, -30, 119, 73, 7, 23, 64, -6, 25, -128, -37, -30, -42, -90, -110, 55, -7, -67, -71, 19, -6, 66, 103, 110, -120, -21, -89, 25, -126, -75, 98, -128, 23, 89, 73, -98, -16, 10, 24, -118, 10, 115, -20, 97, -102, -2, 24, 19, 59, 81, -90, -75, 19, -115, -92, 27, -7, -53, -76, -5, 0, -106, -5, -105, 111, -59, -74, -32, 79, 78, -22, -39, 66, 86, -70, 92, -43, 82, -17, -112, 35, 22, -58, -74, 35, -22, 81, -100, 53, -123, 24, -74, -101, -109, -51, -117, -40, 3, -21, -89, -46, 85, 1, -108, 43, 59, 112, -128, 14, -33, -111, -79, 117, -41, -24, 25, 65, -71, 53, -10, -65, -51, 44, -38, -31, 122, -27, 57, -3, 80, 97, 79, 37, -30, 99, -47, -99, 83, -47, 43, -77, -30, 93, -88, 57, -59, 65, -6, -2, -9, 113, 61, 68, 29, -104, -91, 23, -3, 95, -107, -50, 64, 100, 115, -94, 72, -60, -65, 27, 22, 107, 78, 120, 72, 119, 50, -115, 56, -84, 11, -81, -99, -55, 116, 59, -31, -103, -46, 94, 120, -25, -84, 56, -52, -96, 90, -108, -28, -102, 47, 122, -123, -2, 115, 77, -11, 37, 90, -83, 81, -27, -35, 111, 46, -47, 42, -113, -22, 124, 110, -29, -28, -102, -101, 48, -70, 118, 68, 31, -112, -13, 25, -107, 113, 12, 98, -26, -79, 60, 20, -125, -95, 113, 114, 80, -62, 28, 95, 44, 24, 77, -113, 124, 104, -85, 44, -94, -95, -16, 65, -79, 100, -37, -58, 85, 103, -88, -68, -103, 100, 80, -100, -123, 65, -114, 85, -125, 42, 53, 47, -62, 2, 63, -65, -22, 106, 107, 13, -117, -36, -50, -68, -64, 41, 2, -107, 17, 42, -47, 42, 14, -95, 70, 19, 98, 84, -23, 101, -2, -98, 21, 64, 32, -44, 127, -117, -66, 107, 24, -55, -57, 102, 5, 7, 16, -121, 28, -95, 49, 110, 75, -65, -113, 17, 82, 114, -27, -69, 87, 99, -39, -20, 35, 122, 64, 35, -123, 126, 14, 29, -57, 85, 3, 76, -36, -109, 83, 120, -76, 4, 102, 127, 67, 118, 16, 22, 104, 117, 81, 63, 88, -85, -84, -4, -91, 108, -97, -86, 107, 45, 71, -78, 2, -54, 127, 94, -34, 82, 86, 18, -41, 61, 18, -102, 51, -94, 48, 27, -104, 2, -38, 112, 45, 6, -20, 82, -13, 11, 124, -34, -72, 67, 16, 58, -115, 15, 24, -21, -30, -17, 126, 57, -84, 16, 83, 95, 50, 4, -6, 74, -122, 84, 59, 51, -37, -89, 5, 78, 51, 1, -84, 107, -60, 60, 38, -47, -52, -66, 61, 46, 45, 59, -25, 89, -53, -70, 56, 125, 62, -78, 72, 68, -121, 3, -9, -30, 42, 124, -80, -35, -3, -36, -55, 65, -104, 111, -109, -28, -83, 80, -110, 91, 11, -7, 52, 86, 52, -19, 83, -14, 31, 27, -73, 38, -98, 46, -120, 73, 43, -72, -90, -88, 20, -17, 106, 45, -34, 125, -111, 12, 77, -92, -25, -40, 29, -101, -82, -47, 8, -127, 68, -88, 29, 123, 78, 59, 41, 87, 4, -44, -113, 43, -3, 36, -102, -25, -47, -7, -28, -30, -123, -79, 6, -20, 9, -92, 7, 55, -11, -112, 56, -71, -72, -43, -76, -122, -111, 94, 93, 21, -78, 109, -64, 47, 17, -37, -106, 98, 84, -6, -60, 89, 43, 75, -59, -76, 111, 76, 107, -28, 92, 36, 30, -108, 121, 82, -101, -118, 48, 120, 32, 99, 101, 96

	
	);

    signal scenario_output : scenario_type :=(-21, 9, 55, 46, -97, 74, 94, -92, -128, 127, -8, -93, 35, 53, 5, -2, 12, 9, 105, -128, -90, 127, -79, -52, 127, 32, -111, 23, -52, -107, 127, -8, -86, 41, 40, 32, -83, -6, -56, -28, 116, -92, 64, 103, -7, -92, -48, 44, -76, 29, 26, 21, -40, -8, -3, -43, 35, 42, 127, -61, -27, 109, -30, -86, -37, 57, -88, 79, 6, -128, 47, 87, -6, -88, 47, -7, -21, 127, -6, -62, -22, 63, -51, -55, 53, -87, 88, 39, -7, 15, 18, -8, -57, -6, 96, -100, -128, 19, 127, 23, -117, -7, 116, 55, -102, -26, 48, 93, -78, -98, 31, 96, -78, -8, 38, -57, 91, 76, 14, -78, -56, 72, -85, -107, 76, -15, -45, 97, -36, 87, 110, -126, -77, 42, 125, -38, 8, 15, -91, -61, 75, 90, -10, 27, -80, -123, 10, 11, -35, -1, 95, 58, 31, 4, -18, -88, -3, 119, -39, -8, 44, -78, -95, -30, -25, 1, 92, 127, 10, -128, -77, 89, 125, -94, -62, 54, -59, 98, 26, -102, 127, -77, 0, 127, -70, 13, -125, -25, 97, 31, -41, -37, -36, 20, 81, -106, 53, 10, -122, 71, 11, -54, 127, -59, -105, 90, -41, 60, -44, -7, 127, -128, -37, 127, 0, -72, -42, 108, -109, -124, 127, 6, -14, 107, -128, -77, 6, 79, 78, -117, -40, 93, 49, -116, 43, 124, -37, -128, 0, 110, 23, -54, 0, 13, -69, 4, 127, -116, -66, 30, -43, 39, 44, -22, -75, 113, 40, -75, 39, -63, 3, 127, 22, -105, -125, 110, -11, 0, 104, -17, -47, -21, -27, -78, 127, 48, -75, 92, -26, -111, -97, 127, 73, -93, 100, 24, -128, -4, -43, 56, 77, -45, 43, -83, 45, 64, -17, 64, -96, -58, 48, 52, -124, 26, 3, -128, 82, 124, -99, 27, 127, -128, 3, 82, -71, 97, -113, 25, 44, -128, 79, 87, 29, -76, -128, 114, -9, -128, 127, 51, -22, 9, -81, 88, -6, -105, 119, 69, -128, 59, 127, -128, 90, 83, -115, 55, -43, 8, 35, -29, 83, -85, -83, 120, -7, -37, 4, -11, 35, -80, 87, 2, -69, 41, -128, 125, 78, -13, -2, -57, 77, -99, -24, 120, -9, -109, -8, -47, 96, -17, -68, 127, -99, -115, 73, 88, 25, -119, -65, 63, -2, -18, 38, 116, -25, -60, 78, -96, -29, 39, 45, 3, -54, 53, -60, -53, 103, 76, -104, 2, 99, -128, -5, 5, -62, 22, 104, -43, -89, 36, -11, 96, -30, 62, 11, -15, 29, -97, -63, -30, 105, 127, -32, -104, -2, 98, 21, -96, 28, -41, -87, 100, -23, 56, 61, -55, -78, -18, 96, -26, 11, -73, -76, -12, 127, 80, -30, -13, -9, 83, -55, -63, 61, -48, -128, 69, 21, 18, 123, 6, 8, -127, -42, 25, -63, -8, 127, 2, -28, 32, 20, -27, -32, -61, -34, 108, 20, -34, -93, 59, 13, 47, -10, -103, 8, -18, 111, 25, -128, 88, 34, 46, -82, 1, 65, -128, 27, -25, 96, -48, 18, 110, -71, -17, 12, 115, -109, -108, 88, -42, 96, 95, -128, -60, -1, 14, 71, 70, 34, -58, -3, -78, -8, 109, -116, 28, 127, -97, -128, 60, 44, 48, -62, 22, 21, -43, 127, -85, -116, -5, 106, -25, -127, 127, 54, -128, -28, 127, -32, -128, 117, 116, -72, -83, 42, 41, -60, -26, 127, -71, 26, 31, -128, 8, 22, 9, 127, -79, -26, 24, -78, 76, -36, 20, -4, 27, 70, -39, 2, 38, -1, -76, -22, 123, -19, 17, -30, -40, 22, -113, 127, 4, -109, 127, -34, -54, -4, -64, 62, 114, -83, 19, -9, -75, 32, -46, 127, 54, -55, -19, -51, -48, 57, 109, -122, -103, 127, 4, 5, 111, -76, -23, -71, 47, 72, -94, -7, 35, 23, 48, -45, -14, 57, -49, -92, 55, 124, -128, -30, 76, -13, 63, 21, -110, -10, 90, -34, -73, -49, 14, 5, 35, 127, -71, -70, 25, 29, 62, 55, -104, -34, 9, 77, -19, -34, 14, -128, 102, 17, 8, -56, 51, 62, -28, -65, 58, 55, -93, -17, -26, 110, -59, 43, 46, -87, -36, 79, -62, 32, 127, -128, -5, 127, -91, -20, 109, -110, 57, -26, -44, 55, -77, 5, 87, 76, -71, -12, -12, -128, 127, 105, -55, -90, 3, -1, -18, 117, 32, -51, -7, -24, 17, -20, -102, 127, -51, -128, 60, 127, -52, 13, 23, -89, 45, -72, -1, 127, 63, -59, 6, 29, -100, -42, 97, 48, -49, -79, 15, 22, -128, 20, -29, 52, 127, -128, 20, 96, -87, -115, 77, 90, -111, -77, 9, 93, -4, 2, 69, -91, -17, 80, -93, 78, 32, -128, 127, 127, -70, -36, -23, 36, -64, -42, 86, 44, 44, -93, 0, -40, -11, 37, 21, 63, -90, 69, -42, -51, 64, -6, 42, 41, -122, -6, 114, -125, 40, 52, -128, 14, -20, 42, 6, -74, -6, 99, -36, 44, 0, -30, -1, -5, 0, 25, 52, -82, 89, 9, -103, -32, 47, -54, -19, 85, 127, -128, 8, 127, -85, -89, -48, 96, 95, -47, -128, -57, 54, 22, -53, 26, 127, -65, -128, -7, 127, 59, -97, 90, -117, 35, 11, -96, 127, -17, -128, 103, 73, -128, 81, 0, -97, 127, 88, -128, -53, 127, -72, 0, -25, -81, 19, 117, 40, -128, 127, -4, -63, 81, -128, 56, 66, -120, -2, 9, 58, 14, -116, 127, 31, -78, 127, -37, -59, 36, 36, -123, 3, -25, 34, 123, -113, -100, 57, 117, -83, 6, -31, -103, 56, -9, 104, 79, -93, -95, 94, 127, -128, 13, 91, -56, -37, 38, -48, -94, 85, -44, -15, 42, -60, 15, 127, 8, -94, 37, -60, 55, 0, -121, 127, 7, -94, 47, 93, -7, -57, 35, -46, 43, 39, -128, 30, 8, -128, 127, 59, -46, -92, 48, 127, -128, -89, 126, 37, 0, -70, 24, 45, -68, -60, -35, 127, 24, -128, 89, 18, -44, 79, -22, 29, -69, -114, 30, 97, -59, -17, -21, 85, 69, -128, 81, 98, -74, 10, -8, -34, -53, -11, 127, 24, -79, -20, 15, -52, -6, 60, -27, -19, -45, -1, -21, 47, 34, -30, 127, -30, -58, 127, -108, -128, -11, 127, 110, -93, -10, -82, 68, 77, -102, 83, -46, -128, 31, 127, -43, 23, -3, -25, -2, -81, 127, -73, 0, -5, -58, 127, -34, -82, 59, 58, -75, 41, 30, -111, -45, 127, -9, -128, 73, 83, 61, -18, -21, -69, -36, -19, -77, 122, 99, -87, -114, 76, 37, 31, 26, 12, -35, 34, -41, -128, 104, 40, 30, 91, -38, -128, 81, 127, -128, -41, 81, -60, -53, 32, 32, 58, -30, -11, 22, -114, 96, 49, -43, -25, -63, -9, 127, 85, -128, -79, 121, 76, -44, -5, 21, -80, 17, 63, 35, 38, 15, -80, 23, -47, -40, 49, 17, -78, 43, 34, -128, 127, 52, -42, 68, -17, -24, 51, -116, 2, 113, -1, -78, -76, 0, 102, -11, 9, 6, -127, 94, -11, -7, 73, -53, -17, -60, -28, 100, -57, -21, 103, 30, 61, -103, -49, 85, -122, -26, 127, 63, -109, -13, -7, -31, 127, -128, 3, 127, -128, -89, 39, 90, -107, -65, 47, 35, 18, 15, -56, -31, 127, 35, -128, 91, -64, -11, 127, -128, -2, 37, 83, 29, 15, -82, -128, 127, -30, -128, 127, 32, -55, -7, -55, 34, 71, -47, 66, 79, -3, -128, -98, 127, 37, -69, 32, 15, -51, -55, 36, 87, -23, -38, -28, -1, 32, 10, -45, 45, -107, -85, 90, -4, 52, 27, -125, -63, 127, -68, -128, 127, -64, -74, 127, 15, -116, 8, 38, 24, -52, -105, 117, 114, -128, -90, 119, 76, -86, -106, 127, -39, -3, -11, 4, 42, -14, 63, -27, 2, -2, 29, -18, -23, -15, -43, -1, 57, -39, -128, 93, 61, -62, 18, -2, -19, 107, -79, -85, 23, 10, 3, -4, 0, 0, -5, 48, -22, 63, 14, -17, 92, -128, 11, 34, 40, -75, 42, 96, -128, 127, -48, -41, 54, -23, -49, 40, 76, -123, -45, 70, 75, -86, 62, 70, -97, 88, -79, -75, 127, -62, -57, 12, -3, 95, 44, -128, 63, 76, -60, -51, -17, 91, 48, 29, -91, -128, 76, 127, -124, 28, 17, -8, -28, -103, 66, 70, -58, -2, -7, 51, 120, -76, -94, -29, 25, 103, -6, -106, 38, -64, 38, -23, 37, 80, 11, -59, -62, 125, -128, 51, 106, -113, 39, 41, 6, -92, -29, -46, 62, 108, -1, 23, -119, -52, -42, 107, 5, -38, -1, 12, 85, -10, 20, -40, -76, 35, 92, -128, -56, 127, 89, -128, -107, 127, 91, -128, 48, 54, -128, 106, 127, -128, -53, 56, -55, 91, -70, 0, 42, -65, 6, 127, -45, -128, 99, 30, 68, -42, -65, 38, -78, 34, 45, -2, -26, -46, 86, -21, -23, 122, -112, -39, 127, -24, 9, -46, -116, 127, 94, -79, -89, -43, 56, 18, -11, -78, 98, 45, -114, 30, 53, -5, 20, 93, 18, -128, -99, 110, -36, 63, -2, -99, 19, 124, 97, -128, -69, 21, -28, -2, 105, 26, -48, -31, 52, 119, -116, -41, 127, -49, -17, 26, -15, 30, -63, 12, 17, 24, -110, 29, 78, -106, -76, 104, 14, -10, 121, -98, 8, 80, -73, -44, -76, 73, 64, -26, -4, -9, -40, -21, -12, -89, 127, 116, -63, -53, -20, -3, -63, 69, -13, -11, 127, -100, -68, 12, -66, 15, 110, -63, -82, 46, 45, 25, -76, -30, 4, 77, 108, -75, 53, 85, -128, 59, 51, -128, 12, 3, -2, 98, 27, 15, -76, 28, -82, 52, -2, -128, 66, 75, -13, -58, 120, 24, -39, 38, -15, -7, -46, -57, -43, 12, -4, 19, 32, 19, 45, -1, 54, -119, -53, 123, -100, -119, 121, 15, -107, 91, 62, -45, -25, 48, 112, -105, -71, 112, -65, -77, 77, 49, 10, 31, -128, 51, 41, -94, 63, 89, -64, -64, -23, 79, 17, -128, 127, 89, -103, -117, -3, 127, -21, -35, 51, -96, 93, -69, 26, 21, -128, 102, 34, 97, -103, -51, 127, -59, -112, 18, 39, -19, 98, 9, -94, -72, 93, 4, 27, -15, -106, 21, 107, 56, -19, -37, 3, 63, -99, 27, 48, -17, -70, -58, 82, 18, -115, 40, -35, -30, 17, -22, 127, 66, 19, -120, -128, 119, 43, 26, 58, -31, -114, 15, 63, -128, -10, 40, 90, 73, -127, -2, 57, -4, -68, -39, 19, 12, -38, -42, 127, -70, -34, 127, -128, -7, 127, -115, -85, 76, -49, -20, 13, 36, -44, 51, 87, -64, -66, 30, 9, 2, -15, 78, -8, -77, 37, -20, 125, -49, -27, 95, -80, -29, 13, 5, -44, -23, 90, 15, 12, 32, 22, -128, -75, -14, 72, 127, -87, -128, 6, 120, -4, -10, 1, 30, -98, 41, 41, -128, 39, -18, 96, 106, -53, -46, -34, -95, 124, 11, -73, 127, -128, -1, 1, -58, 127, -121, -41, 87, -115, 127, -27, -71, 127, -19, -46, 37, 15, 1, -125, 24, 127, -39, -27, -36, -43, -97, 69, 36, -78, 30, -19, 18, -13, -44, 127, 104, -128, -53, 3, -14, 51, -18, -54, -2, -30, 94, -8, -3, 90, -128, 52, 70, -128, 30, 5, -9, 83, 34, 19, 37, -128, 44, 44, -128, 30, 8, -31, 55, 103, -35, -114, -29, 127, -23, -73, 110, 60, -55, -52, -37, 45, -43, 4, 104, -57, 9, 82, 54, -119, -42, 94, -60, 0, -78, -7, 127, -112, -4, 31, 32, -49, -75, 0, 61, 83, -82, 17, -39, 57, 107, -78, -93, 103, -46, -128, 56, 117, 93, -85, -128, 94, -26, -6, 49, -98, 20, 1, 26, -30, 44, 53, -75, -37, 60, -14, 13, 127, -45, 6, 59, -89, -30, -26, -12, 85, -55, 37, 43, -108, -44, 93, -57, -62, 83, -38, 26, 60, -39, 42, 57, -128, -88, 127, -44, -68, 127, -3, -65, -37, 43, -3, -115, -14, 127, 55, -127, -69, 98, 75, -30, 49, -27, -43, -18, 24, 100, -1, -72, -88, 85, -46, -78, 127, 87, -92, -81, 95, -55, -128, 28, 127, 1, -93, -18, -55, 127, -3, -126, 63, 74, 59, -86, -94, 22, 49, 113, -73, -92, 42, 35, -47, -35, 127, -100, -90, 88, 12, -35, 5, 56, -11, -36, 63, 74, -64, -128, 47, 124, -91, -83, 55, -24, -10, 107, -8, -115, 37, 114, -66, 78, -46, -74, 73, -90, 26, 126, -8, -119, -55, 2, 95, 78, -39, 1, 6, -103, 53, 10, 30, -44, -65, 79, -68, -41, -34, 124, -15, 0, 41, -37, 68, -3, -76, -78, 106, 91, 43, -98, 17, -21, -89, 107, 58, -97, -74, 71, -4, -65, 93, 19, -104, 24, 68, 15, -65, 70, -60, -37, 63, -49, 112, 83, -18, -128, 48, 77, -65, 87, -13, -54, 65, -73, -128, 127, -17, -17, -23, -10, 100, 21, 39, -128, -99, 115, 2, 22, -45, -47, 127, -28, -66, 119, -91, -82, 127, -87, 1, 117, -128, 31, 69, -128, 122, 83, -20, -54, -83, -2, -63, 26, -9, 127, 5, -111, 61, 14, 90, 5, -128, 75, 127, -72, -2, -68, -110, 113, 40, -110, 12, 52, 66, 38, -64, 26, -27, -41, -58, 52, 100, -125, -117, 127, 3, -105, 21, 28, 127, -85, -128, 127, -19, -128, 113, 127, -81, 1, 53, -1, -80, -121, 95, -11, -76, 40, -11, 58, 127, -78, -43, 61, -9, 18, 0, -128, -80, 127, 64, -128, -91, 127, -12, -100, -13, 107, 29, -94, 127, -104, -46, 22, -25, 7, -14, 85, 0, 3, -14, -38, 119, 121, -128, -32, 127, -18, 1, -128, 15, 72, -117, 113, -9, -82, 2, -18, 22, -3, 112, -75, -59, 58, -83, 103, 18, -63, -8, 25, 120, -34, -128, 92, 88, -128, 51, 49, -122, 21, 80, 44, 49, -5, -3, -110, -43, -32, 32, 124, -38, -45, 54, 80, 2, -128, 37, 24, -54, -15, 61, 62, -87, 112, -46, -128, -31, 127, 56, -128, -7, 127, 106, -128, -8, 104, -72, -96, 80, -45, 32, 36, -89, 119, -66, -78, 127, -73, -42, 65, -83, 15, 92, 55, -105, 56, 95, -128, 64, -36, -70, 9, 113, 27, -128, 104, 100, -30, 0, -13, -31, 22, 23, -89, -41, -36, 28, 41, -100, -15, 76, 0, -6, -23, 61, 68, 26, -39, -36, 81, -69, -114, 97, 38, -83, -12, -41, 23, 127, -47, -128, 126, 127, 37, -128, -54, 6, 27, 127, -128, 47, 11, -93, 30, -4, -38, 104, 14, -74, 99, -86, -128, 127, 127, -102, -94, -38, 48, 113, -122, 10, 123, -5, -14, -26, 69, -117, -13, 127, -128, -103, 127, 5, -45, 127, -5, -57, 76, -128, -88, 127, -66, -37, 94, -88, 57, 127, -128, -46, 66, -24, -46, 9, -24, 127, -23, -128, 60, -69, 127, 37, -128, 105, 45, -3, 39, -106, -15, 85, -87, 82, -5, -106, 39, 53, 26, -98, 14, 85, 34, -109, -119, 127, 42, -128, 122, 20, -62, -54, 0, 83, -53, 51, -49, 40, 37, -3, -71, 26, 74, -128, 108, 31, -36, -52, -55, -2, 7, 106, 79, -128, 2, 127, 21, -113, -128, 127, 65, -69, 89, -92, -128, 42, 111, 2, -112, 6, 1, 12, -5, 44, 82, -97, -64, 52, 8, 29, 3, 47, -21, -104, 127, -29, -128, 127, 10, -107, 79, 83, 45, -69, 38, -96, -20, 127, -86, -128, 121, 97, -128, -38, -41, 127, 5, -107, 5, 20, 103, 0, -85, -103, 90, 127, -128, -17, 127, -125, -97, 43, -30, 106, 124, -36, 41, -59, -36, -42, 1, 40, 65, -128, 7, 18, 13, 7, -81, 12, 35, 18, -20, 127, -94, -83, 127, -40, -107, 63, 34, -59, 62, 35, -115, 37, 39, -72, -10, -29, 85, -53, 20, 127, -128, 22, 127, -128, 36, 80, -128, 68, 64, 47, -36, 13, -8, -85, -20, 80, -65, 23, 13, 3, 53, -95, 39, 60, 15, 17, -124, -87, 127, -112, -122, 14, 106, 3, -128, 127, 47, -86, 7, -28, -31, 127, 127, -46, -113, -36, 35, 17, -56, 60, 14, 2, -40, 56, 95, -128, 85, 125, -107, 48, 22, -49, 58, -62, -44, 125, -123, -128, 44, 43, -20, 5, 20, -74, 127, 48, -112, 0, 68, 48, -128, -57, 53, 13, -40, 116, 26, -128, 58, 127, -112, -97, 110, 99, 22, -126, 44, 92, -85, -103, -42, 90, 48, -66, 52, 2, 26, -70, 7, 93, -53, 49, 25, -128, -120, 127, 104, -98, -128, 15, 56, -82, 64, 127, -128, -61, 74, -91, 3, 127, -47, -41, 48, 2, 109, -98, -128, 127, 22, -128, 47, 13, -77, 45, 18, -12, 36, -56, 83, 48, -41, -54, 5, 55, -115, 63, 127, -86, 3, -13, -119, 127, 85, -75, 0, 5, 55, -128, -35, 85, -85, -27, 72, 25, -25, 88, 5, 0, 59, -73, -97, 24, 29, 57, 36, -54, -41, 26, -96, -69, 127, -31, -110, 71, 123, -120, -102, 127, -74, -128, 52, 40, -21, 83, 59, -19, 9, -85, 22, 34, 37, -81, -125, 112, -22, -77, 29, 98, 94, -72, -126, 80, 88, -55, -38, 26, 54, -128, -5, 127, -128, 43, 24, -123, 117, 86, -112, -59, 45, -87, -14, 55, -5, 9, 127, -34, -40, -4, -81, 59, 76, -23, -54, 22, -76, 103, 8, -49, 127, -7, -27, -128, 42, 127, -91, -30, 53, 26, -98, -119, 127, 27, -64, -61, 81, 52, -89, 39, 10, 49, -100, -53, 32, 2, 115, -45, -92, 127, -69, -128, 127, 56, -106, 18, 23, 31, -23, -104, 69, 32, -34, -19, 70, 79, -91, -5, -18, -128, 1, 127, 58, -102, -90, 98, 79, 14, -106, -128, 127, -20, -107, 123, 42, 4, -59, -75, 42, 71, 4, -85, -37, -26, 88, 25, -128, 44, -10, 12, 53, -14, 14, -71, 75, 104, -128, 12, 126, -121, 42, 77, -97, -36, 12, -6, -63, 116, 62, -27, 29, -81, -66, -43, 91, -19, -44, 127, -23, -19, -38, 74, -45, -21, 34, -128, 93, 19, 46, -13, -53, 83, 30, 31, 36, -114, -124, 17, -28, 103, 127, -5, -128, -116, 127, 99, -128, -51, 64, 29, 70, 19, -53, -121, 3, 127, -87, -128, 127, 127, -128, -45, 73, -87, -7, 81, -38, 18, 54, -36, -41, 43, -35, -20, 111, -80, -100, 127, 7, -42, 38, -71, 20, -51, 8, -15, 56, 105, -128, 68, 55, -83, -22, 100, 11, -36, -12, 13, 9, -128, -10, 127, 47, -53, -48, -24, 58, 30, -54, -74, -5, 127, 4, -24, 88, 2, -12, -17, -42, -128, 56, -19, -19, 28, -97, 3, 127, 73, -128, -22, 124, -6, -88, -6, 127, 3, -38, 41, -128, 103, 108, -128, 86, -37, -128, 127, -27, -128, 127, 87, -92, -41, 79, 72, -57, -23, 103, -69, -128, 124, 49, -11, -78, 1, 7, -126, 17, 127, 61, -128, 77, -17, -64, 120, -87, 14, 61, -108, 90, -44, 27, -11, -80, 100, 60, -106, -106, 127, -20, -56, 102, -115, -23, -9, 47, 127, -128, -89, 74, 112, -42, -78, 100, 109, -128, -126, 127, 56, -45, -11, 59, -28, -19, -26, 78, 34, -128, 7, -12, 44, 127, -128, -21, 99, -128, 62, 8, -94, 117, 42, 15, 63, -7, -40, -9, 24, 10, -74, -63, 4, -80, -31, 127, 44, -64, 63, -108, 39, 22, -114, 121, -68, -22, 55, 4, 10, 72, 6, -55, 27, -99, 1, 94, -100, -34, 91, -64, -48, 127, 21, -83, 92, 17, -108, -12, -2, -80, 79, -2, -86, 127, 70, -119, -66, 127, 65, -65, 44, -76, -76, 41, -17, 112, -96, -69, 71, -37, 48, 11, -17, -79, -26, 42, 99, 9, 27, -98, -26, 102, -128, 113, 15, -19, -14, -43, 105, 52, -77, -32, -17, 41, -35, -24, 127, -128, -59, -1, 31, 127, 4, -128, -128, 127, 44, -37, 28, -114, 96, -41, -43, 127, -128, -128, 127, 7, -28, 76, -85, -61, 11, 59, 126, -28, -119, 90, 35, -36, 82, -90, -49, 93, -75, 4, 31, 14, -5, -127, -51, 60, -10, 93, 10, -128, 108, 127, -90, -78, 24, 20, 0, 29, -77, -19, 2, 0, 26, 45, -4, -73, -34, 103, 127, -115, -49, 47, -56, -87, 82, 42, -71, 107, -63, -14, -34, 51, 109, -123, 3, -49, -91, 127, 126, -128, -47, 127, 7, -25, -11, 8, 79, -56, -45, 94, -128, -89, 114, -29, 10, -32, 19, 127, -128, 4, 127, -128, 91, 19, -81, 49, -61, 52, -20, 75, 60, -78, 52, -81, -64, 42, -62, -11, 127, 79, -128, 61, -20, -31, 29, -39, 119, 43, -74, -5, 75, -126, -128, 127, 52, -48, -48, 39, -7, -63, 108, 54, -106, -61, 127, -23, -58, 104, -9, -72, -3, 73, -59, -12, 35, -27, -21, -28, 21, 95, -41, -82, -23, 0, 11, 0, 127, -43, -128, 127, 72, -49, -9, 7, -83, -21, -10, 53, 38, -9, -25, 41, 57, -82, 59, -91, -100, 127, 24, -80, 96, 22, -128, -110, 32, 29, 78, -62, -3, 105, 59, -88, -90, 56, 77, -24, -8, 97, -128, -115, 90, 31, -75, -69, 127, 125, -128, -105, 127, 49, -5, 42, -106, 54, 74, -78, -70, -31, 55, 69, 71, -80, 24, -28, -18, 95, -51, 7, -31, 48, -117, -121, 92, -40, -2, 11, 96, 9, -99, 38, 100, -78, -102, 4, 127, 116, -79, -92, -60, -22, 127, -32, -93, 127, -60, -79, 98, -68, -70, 76, -45, -25, 106, 2, -29, -96, 58, 55, -80, -46, 100, 17, -128, 127, 11, -128, 115, 127, -124, 9, 127, -128, 17, 75, -128, 5, -36, 111, 85, -108, -4, 40, 83, -98, -98, 56, 0, -79, 85, 103, -128, -6, 122, -68, -59, 127, -26, -128, 89, 41, 54, -2, -61, 64, 36, 9, -128, -128, 127, 108, -64, -72, 6, 24, -12, 58, 40, -19, 6, -32, -100, 70, 106, -22, 32, -115, -27, 8, -60, 17, 60, -12, 14, 29, -128, 100, 8, -107, 127, -59, -128, 85, 25, 15, 65, 44, -87, -43, 68, -111, 86, 112, -47, 32, -59, 25, -80, -77, 6, 21, 90, 23, 40, -52, -128, 127, 0, -119, 66, -77, 22, 71, -32, 41, 115, -128, -59, 34, -15, 127, -82, -85, 78, 98, -61, -128, 127, 14, -87, 98, 68, -128, -23, 115, -58, 28, 20, -9, -95, 56, 96, -79, -68, 104, -5, -128, 127, 75, -128, 3, 45, -37, 98, -70, -79, 39, -35, 14, 23, 99, -82, -87, 127, 34, 21, -80, -81, 48, 62, 5, -87, -19, 119, 27, -128, 117, 71, -128, 13, 122, -22, 54, -73, -70, -10, 5, 120, -90, 57, -54, 14, 127, -128, -6, 41, -123, 70, 106, -76, -58, 119, 14, -85, 44, 45, -11, -34, -65, 48, -29, -124, 36, 127, -46, -73, 127, -13, -116, -69, 44, 22, -56, -18, 71, 82, -19, -20, -5, -97, 94, 115, -128, -30, 32, 65, -29, 29, 25, -89, 77, -35, -29, 108, -48, -37, 62, -65, -41, 104, 9, 1, -69, -2, -27, 7, 74, -41, -14, 32, 82, -116, -30, 103, -6, 0, -26, 7, 20, 0, -49, -86, -28, 116, -21, -66, 77, 8, 49, 25, -44, -86, 29, 82, -128, 11, 83, -52, -35, 70, 12, -128, -35, 127, 112, -48, -15, -64, 0, 9, -92, 112, 70, -123, 36, 49, 26, -87, -86, 121, -96, 70, -9, -56, 127, -128, -7, 7, 4, 127, -128, 28, 127, -128, 14, 108, -17, -10, -128, -7, 127, -44, -88, 40, 61, -61, -89, 99, 6, 12, -12, -41, 71, -20, -61, -4, 39, 71, -2, -109, 23, 75, -87, -13, 111, -81, -86, 105, 60, -38, -94, 35, 109, -2, -116, -8, 127, -25, -105, -6, -6, 39, 95, 58, -128, -112, 56, 96, -80, 26, 127, -66, -56, -66, -37, 23, 12, 22, 127, -122, 27, 21, -80, 127, -15, 24, -74, -29, 4, -20, 108, -8, -128, 58, 55, -121, 96, 73, -30, 43, -63, -10, 15, -113, -106, 127, 56, -98, 9, -4, 13, -8, 22, -35, -58, 15, 127, 12, -15, -43, 36, 80, -49, -70, -43, 10, 4, 7, 91, 5, -128, 76, -37, 41, 108, -128, 29, -19, -51, 127, -68, -1, -19, -39, 127, -126, 12, 94, -69, -12, 52, 0, -116, 12, 87, -14, 19, -65, -128, 115, 93, -102, -41, 105, -66, 34, 127, -46, -128, -57, 127, -14, -104, 127, -22, -128, 49, -41, 112, 126, -61, 10, -61, 52, 13, -128, 86, 0, -61, 82, 76, 24, 7, -127, -19, -18, -87, 93, 97, -85, 32, 42, -60, -38, -51, 116, -37, -45, 107, -87, -64, 51, 78, 57, -88, -91, 127, -49, -79, 63, 35, 28, -94, 49, 97, -128, 42, 3, -59, 127, -78, 4, -6, -128, 125, 87, -18, -70, -105, 95, 1, -23, 127, -78, -112, 55, 25, -19, -21, 127, 32, -128, -24, 127, 92, -128, 21, 125, -128, -1, 32, 3, -40, -5, 96, -114, -59, 85, -26, -13, 127, -31, -6, 80, -71, -88, -86, 127, 31, -109, 92, 68, -32, -128, 58, 61, -104, 78, -35, -21, 28, 7, -24, -5, 0, 39, 62, -64, -66, 37, 127, -127, -128, 127, 111, -58, 3, 57, -64, -113, -11, 32, -71, 117, 44, -14, -15, -13, 52, -49, -3, -103, -31, 127, 37, -36, 11, -45, -100, 127, -9, -128, 127, -4, -44, 124, -22, -12, -5, -43, -120, -44, 127, -7, -124, 51, -20, 54, -6, 41, 1, -41, 123, -40, -70, 14, -70, 98, 115, -128, 43, 108, -128, 13, 127, -128, -44, 127, 29, -53, -128, 111, 42, 13, -92, -36, 54, -107, 14, 15, 123, -30, 9, 44, -30, -27, -128, 127, 22, -44, -4, -117, 74, 18, 85, -12, -81, 29, 125, -57, -20, 25, -128, 71, 4, -26, -6, 31, 54, -40, 85, -23, -31, 123, -128, -14, 58, -128, 81, 54, 10, 32, -64, 75, 79, -128, -82, 0, 82, -2, -46, 60, -8, 6, 87, -10, 6, -82, -124, 66, 35, 107, 37, -128, 44, 66, -19, 60, -34, -100, -30, -15, 87, 87, -128, 24, -48, -61, 127, -9, -32, -35, -94, -36, 127, 127, -53, -17, -128, 56, 1, -87, 127, 3, -15, 5, -75, 3, 68, -103, -86, 8, 43, 127, 51, -57, -24, 41, -91, -34, 42, 32, 75, -58, -128, 59, 80, -17, -1, -41, 32, 1, -97, 8, 11, 81, -28, -52, 82, 7, 31, -52, 47, -86, -46, 100, 48, -77, -40, 1, -110, 11, 7, 127, 99, -128, 29, 29, -128, -3, 127, 44, -7, -106, -90, 9, 127, 25, -49, 59, -115, 22, 13, -95, 98, 113, 0, -9, -110, -34, 127, -75, -27, -1, -92, 73, 35, -103, 75, 86, -117, 68, -13, -120, 121, 40, -111, 59, 107, -128, -103, 127, 34, -94, -61, -11, 20, 127, -66, -78, 98, 46, 66, -128, -95, -19, 102, 85, -128, 23, -15, -10, 46, -58, 57, 124, -24, -25, 24, -100, 37, 102, -105, -70, 12, -7, 62, 30, -69, 40, -58, 35, 81, 13, -102, -7, -9, 6, 70, -128, 28, 22, 44, 26, -4, -58, 1, 10, -78, -4, 107, -48, -82, 11, 39, 76, -2, -49, -76, 124, 127, -128, 0, 68, -123, 95, 14, -123, 99, 51, -32, -72, -69, 17, 114, 72, -46, -38, -100, 70, 102, -32, 19, 7, 5, -102, -60, 8, 5, 8, 127, -57, -86, 125, -25, 15, -13, -3, 110, -114, -94, 83, -27, -18, 95, -72, -91, 55, 46, -44, 123, -46, -34, 127, -31, -34, 36, -98, -19, 35, -82, 110, -58, 55, -3, -35, 60, -15, -3, -49, 70, 42, 27, -116, -121, 127, -30, -61, 127, 9, -75, 68, 2, -81, 15, -23, 79, 7, -112, 58, 6, 29, -69, -1, 75, -68, -39, 106, 100, -54, -103, 20, 32, -105, 65, 61, -14, 28, 26, -31, -111, -3, 2, 54, 64, -25, 62, -18, -128, -4, 8, 2, 127, -68, -128, 62, 56, -13, -23, -22, 127, 14, -3, -35, -44, 51, 27, -28, -103, 66, 96, -63, 19, 127, -128, -61, 108, 85, -124, -48, 74, -113, -10, 23, 19, -19, 46, 74, -39, 12, 83, -112, 73, 68, -128, 21, 125, -119, -1, 14, -45, 89, -46, 9, -5, 13, -61, -77, 109, -26, 23, 127, -128, 6, 127, -128, 19, 6, -15, -29, 24, 60, -128, 95, 92, -55, -78, 34, 59, -128, 59, 7, -32, 5, 24, -41, -11, 127, -124, -94, 125, 82, 0, 13, -73, 11, -79, -46, -9, 65, 68, 12, -68, -27, 127, -128, -35, 22, 71, -19, -95, 124, -5, -128, 127, 12, -128, 123, 127, -110, 18, 95, -128, 62, 73, -48, 29, 4, -103, 26, 64, -27, 34, -2, -20, -54, 72, -104, -21, 127, -122, -80, 40, 69, -31, -52, 92, -21, 64, 23, -88, 76, 82, -43, -60, 10, -52, -23, -15, 45, -40, 58, 9, 0, 49, -7, -18, -98, 89, 105, -5, -1, -128, -110, 73, -10, -12, 122, -1, -107, -36, 107, 111, 39, -94, -95, 56, 11, 26, 37, -128, 29, 86, -122, 27, 104, 53, -1, -128, -3, 106, 36, -48, -20, -75, -6, 127, -98, -38, -32, -9, 65, 68, -57, -40, -23, 43, -27, 0, 68, -26, 80, -97, -120, 127, 70, -22, 49, -80, -128, 48, 31, -88, -26, 127, -18, -35, 127, -73, -85, 104, -90, -12, 127, -128, -55, 110, 87, -94, -48, 5, -76, 0, 64, -11, -40, -9, 9, -21, 73, 23, -11, 104, -74, -8, 77, -52, -15, 19, -81, -95, 96, -12, 79, 27, -109, 51, -44, -11, 115, 51, -12, -119, -93, 58, 26, 14, 8, 30, 25, -120, 99, 2, -9, 19, 0, 60, -30, 20, -128, 87, 66, -51, -79, -37, 127, -47, 10, -66, -15, 116, -8, -36, 4, -109, 27, 24, -87, 35, 24, 122, -90, -72, 127, -111, -46, 127, -47, -42, -41, 49, -4, 35, -6, -81, 28, -20, -80, 8, 70, 86, -71, -80, 56, 87, -5, -107, -66, 103, 69, -44, 28, 18, -86, -22, 104, 46, -54, -85, 4, 96, -41, -128, 127, 106, -76, -21, -93, 38, 127, -25, -66, 63, 73, -20, -7, -77, -126, 122, -18, -46, 70, 17, -34, -11, 25, -113, 43, 126, -13, -128, 41, 127, -128, -8, 58, 17, -78, -24, 48, 56, -56, -15, 127, -128, 10, 108, -52, -116, 12, 126, 14, -113, 1, -14, 70, -17, -119, 112, 76, 49, -40, -35, 0, 47, -54, -121, 75, 20, 38, -72, -70, 21, -81, 54, 9, 116, -66, -30, 127, -64, -58, 6, 56, -106, 2, 120, -121, -83, 44, 0, -26, -22, 122, 127, -128, -75, 41, 59, 127, -115, -128, 64, 64, -87, 79, 73, 19, 40, -121, 48, 15, -128, 66, 40, -85, 28, 127, -22, -60, -12, -17, 92, -46, -49, 64, -20, 15, 100, -121, 0, -12, -79, 24, 23, 18, 94, -61, -108, 127, 9, -60, -64, 31, 127, -68, -19, 18, -79, -36, 116, 53, -55, 11, 45, -77, -107, 31, 127, -51, -77, 127, -96, 30, 108, -40, -109, 19, 89, -38, -35, -79, 96, 40, -48, 52, 17, -76, 38, 121, -123, 0, -12, 52, 2, -128, -14, 53, 35, 80, -4, -10, 12, -60, 46, -61, -91, 96, 103, -7, -95, -116, 109, 127, -82, -98, 48, -62, 21, 47, 26, 121, -128, -128, 127, 8, -125, 125, 55, -61, 42, -98, -27, 20, 40, -20, -69, 127, 65, -125, -19, -28, -48, 88, -104, 69, 127, -98, 41, -43, -10, 100, -128, 71, -38, -128, 86, 29, -28, -41, 15, -17, 22, 127, -4, -91, -74, 127, -5, 1, 30, -17, -32, -10, 64, -128, 93, -26, 4, 87, -63, 28, -38, 25, 52, -70, -86, -82, 127, 29, -128, 127, 1, -111, 112, 3, -22, 30, -30, 17, 21, 5, -6, -9, 25, -128, -96, 88, 0, 96, -59, -14, 115, -96, 42, -15, -128, 114, 46, 1, -52, -74, 127, -47, -128, 54, 127, 7, -111, -24, 63, -87, -11, 62, -86, -12, 94, -32, 29, 127, -128, 13, 104, -19, -48, -37, -28, -8, 32, 26, -12, -15, -9, -69, 127, -18, -21, 127, -128, -88, 72, 65, -24, 20, 122, -83, -128, 32, 75, 62, -71, -18, 106, -128, 10, 24, -28, 127, 8, -128, 8, 2, -11, 127, -73, -34, -24, -51, 62, -21, 10, 95, 37, 12, -45, 13, -69, 0, 3, 15, 55, -64, 34, -64, 18, -2, -29, -12, 92, 127, -128, -90, 127, 31, -128, -45, 3, -11, 53, 26, -36, 58, 112, 27, -91, -79, 48, -2, 64, 46, -128, -24, -11, 48, 60, -32, 43, 19, -18, -21, 0, 0, 68, -26, -108, -72, 85, 45, -125, 127, 62, -128, 31, 27, -98, 98, 94, -54, -61, 12, -5, -9, -55, -7, 31, 10, -46, 83, 23, -60, 56, 26, -27, -60, 9, 22, 15, 55, 62, -80, 31, -63, 19, 14, -27, -46, -69, 76, 51, 52, -106, -96, 47, -2, 45, 40, 1, 29, -76, 70, -40, -13, 90, -65, -42, -83, -36, 127, -35, -128, 96, 127, -34, -79, 25, -56, 30, 102, 13, -76, 8, -89, 23, 12, -81, 68, 21, 108, 48, -22, 14, -128, 6, 70, -6, -79, -6, -7, -128, 127, -21, -39, 113, -15, -88, -82, 127, 85, 12, -15, -128, 26, 53, 37, -4, 3, -57, -128, 127, -5, -128, 127, 49, -128, 25, 48, -26, -20, 11, 26, 93, -14, 19, 5, 12, -78, -71, 127, 7, -21, -107, 109, -43, -43, 127, -46, -4, -128, 58, 97, -128, -49, 10, 107, -47, -2, 127, -86, 6, -34, -13, 90, -46, 37, -88, -23, 111, 23, -85, -21, 3, 4, 42, -34, -6, -4, -31, -46, 52, -12, 23, 96, -111, 71, 3, -115, 61, 121, 20, -128, -55, 12, 112, 80, -128, -116, 63, 124, 52, -27, -55, -89, -15, 127, 22, -25, -51, -2, 111, -46, 15, -27, -99, -52, 11, 66, -21, 66, 28, -128, -57, 127, 11, 53, 17, -89, -74, 87, 27, -14, 57, -59, 79, 29, -71, -43, 6, 70, -53, -65, 66, -35, -82, -60, 75, 78, -38, 89, -49, -2, 121, -117, -27, -17, -20, -41, 54, 49, 39, -74, -110, 98, 58, -37, -49, -5, 110, -48, -115, 68, 43, 100, -6, -44, 68, -95, -115, 74, -41, 29, 64, -104, -38, 4, 40, 86, -39, -99, 127, -10, -128, 69, 56, 77, -15, 37, -87, -89, 127, -61, -27, 71, -111, 4, 32, -70, 72, 66, -40, 62, -60, -128, 127, 42, -128, 3, 127, -18, -104, 125, -22, -89, 127, 64, -128, -15, 109, -107, 81, 61, -120, 46, 96, -9, -128, -51, 116, 71, 8, -78, -49, 127, -59, -87, 4, -21, 60, 99, -44, -9, 23, -27, -72, -12, 43, -48, -71, 125, 27, 4, -9, -52, 79, -97, -51, 94, -2, 59, 6, -128, -17, 127, -41, -65, 62, -68, 96, 113, -126, -94, 105, 93, -128, 44, 73, -116, -11, 8, 2, 22, 6, -1, -31, 54, 85, -89, -47, 127, -39, -34, -17, -51, 111, -52, -120, 127, 63, -28, 58, -22, -95, -19, 77, -70, 22, -65, 12, 127, -63, -128, -8, 127, 1, -46, 40, -96, 56, 127, -128, -126, 127, -28, 10, 24, -74, 109, -34, -128, 125, -11, 22, -13, -21, 93, -78, -4, 28, -29, -73, 127, -26, -85, 109, 13, -99, -76, 127, -49, -121, 127, -34, 20, -38, 21, 32, -107, 127, -37, -36, 14, -1, -25, 6, -23, 36, 111, -40, -89, -106, 120, 27, -122, 32, 105, 76, -76, -125, 44, 65, -62, -2, 79, -54, -34, 95, -18, -106, 1, 127, 0, 14, -53, 17, 11, -74, 86, -64, -65, -38, 29, 13, -37, 91, 37, -86, -15, 127, -30, -128, 38, 97, 15, -115, 92, -29, -13, 68, -128, 23, -12, 104, -9, -55, 116, 4, -95, -19, 127, -19, -60, -20, 0, 81, 64, -128, 35, 75, -128, 13, 69, 0, 72, 78, -83, -35, 93, -105, 1, 127, -91, -128, 64, 91, -41, -10, -83, 55, 127, -128, -106, 95, -5, 77, -14, -125, 127, -24, -76, 127, -58, 23, -9, -128, 105, 98, -128, 18, 0, 22, 119, -85, -111, 0, 15, 4, 127, -73, -93, 98, -14, -54, 127, 10, -128, -54, 121, -27, -72, 79, -100, 108, 55, -105, 6, -23, 3, -8, 127, -1, -128, 76, 105, -68, -128, 127, 116, -31, -98, -123, 73, 39, 10, -6, 60, 56, -66, -14, 68, -107, -128, 127, 127, -108, -90, -35, 64, 55, -45, 13, 55, 30, -110, 19, -35, -68, 108, 91, -102, -22, 127, -38, -128, 12, -5, -73, 42, 85, 99, -119, -15, 127, -128, -15, 58, -85, 97, 79, 2, -111, -56, 102, -116, 34, 77, -128, -35, 127, 127, -128, -23, 102, 4, 19, -114, 9, 126, -81, -59, 37, 28, -81, -22, 116, -128, 45, 25, -45, 127, -128, -109, 69, 100, -41, -89, -1, 12, 15, 127, -51, -87, 115, 53, -49, -53, -15, -34, 40, 98, -99, -100, 127, -27, 63, 18, -126, 99, 46, -128, 34, 82, -64, -89, 3, 89, -31, -38, 94, 17, -90, 83, -42, -128, 127, 61, -23, -102, 75, 10, -34, 127, -100, -55, -13, -29, 117, 43, -123, -19, 127, -98, -115, 81, -28, 38, 125, -28, -128, 74, -9, -56, 119, -83, 9, 29, 25, -24, -64, 94, -11, -63, 31, 87, 22, 10, -100, -5, 55, -31, -26, -24, 70, -1, 49, -117, -108, 127, 7, -83, 22, 42, -108, -79, 127, 42, -52, -11, 58, -89, -100, 57, 0, 114, -51, -119, 127, 39, -128, 3, 19, 0, 125, 82, -128, -8, 127, -82, -22, 19, -126, 5, 32, -71, 77, 127, 3, -128, -8, 69, -69, 39, 81, -31, -41, 31, 65, -111, -107, 127, 34, -94, -25, 12, -9, 11, 2, -70, 127, 126, -95, 38, -68, -17, -43, 14, 125, -38, -91, -68, 36, 31, -34, -60, 9, 80, 122, 32, 2, -128, 19, 38, -44, -46, 24, 127, -78, 21, 89, -112, -3, 34, -71, -60, -14, 80, -52, -70, 53, 14, 10, 49, 44, -28, -15, 44, 78, -56, -68, 82, -11, -54, -57, -47, 57, 113, 77, -128, -11, 127, -98, -17, -13, 29, 63, -30, -81, 17, 78, -38, -125, -55, 18, 78, 60, -3, -34, -10, -21, -95, 44, 127, -3, -19, -77, -96, 127, -35, -75, 87, 103, 46, -128, -56, 116, -64, -80, 42, -36, -29, 127, -14, -88, -10, 107, -38, -7, 65, -43, -35, -23, -4, 99, -32, -15, 15, -124, 120, -55, 21, 5, -93, 75, 28, 37, -37, -24, 127, -39, -68, 127, -73, -39, 41, -77, 61, 9, -92, 127, -38, -123, 104, -37, -28, 76, -56, -44, 127, 14, -64, -34, 26, 25, -3, 54, 53, -13, -128, 8, 127, -18, -45, -80, -12, -40, 40, 8, -60, 127, -96, -52, 45, -23, 98, -27, 49, 31, -45, 27, -98, -104, 127, 73, -83, -9, -22, 12, -59, 43, 14, -100, 35, 127, -31, -18, 87, -1, 17, -128, -9, 117, -43, 29, -64, -95, 41, -12, -53, -30, 127, -5, -128, 127, 69, -3, -72, -95, 10, 64, -91, 0, 127, -65, -29, -32, -44, 57, -23, -54, 81, 127, -128, -104, 127, -43, -9, -2, -45, 115, -44, -21, -77, 48, 106, -128, 92, -1, -87, 64, 31, 43, -128, 38, -15, -8, 127, -62, -128, 127, 62, -66, 87, -29, -128, 51, 123, 30, -128, -64, 127, 0, -92, -110, 58, 127, -114, -79, 127, -21, -24, 55, -128, 72, 44, -128, 99, -25, -41, 127, -126, 70, 62, -32, 32, -73, 49, -27, -36, 93, -99, -66, 104, -37, 6, -28, -47, 83, 71, -66, -78, 52, 127, -59, -68, 3, 0, -12, -48, 127, 78, -128, 52, -7, -128, 54, 81, 61, 19, -112, 9, -77, 15, 70, -105, 21, 7, 29, 99, -116, 6, 10, -58, 127, -46, -94, -36, -36, 47, 97, -82, -53, 127, 111, -65, -128, 13, 56, -72, 6, 106, 83, -77, -30, -32, 52, -59, -19, 120, -128, 102, 78, -128, 79, 0, -13, 127, -81, -12, -18, 22, 82, -81, 12, 48, -128, 68, 19, -79, -9, 28, 57, -114, 0, -9, 52, 7, -58, 30, 91, -22, -62, -9, 5, 127, -15, -128, 105, 93, 3, -110, -25, 90, 0, -13, -82, 92, 5, -53, 5, 1, -27, 30, 75, -76, 56, -73, -23, -11, -36, 64, -65, 89, 5, -24, 51, -8, 30, -44, -56, 37, 37, -88, -52, 47, 51, 47, -55, -85, 0, 107, 61, -32, -18, -12, -64, 1, 114, -128, 0, 72, -65, -35, -21, -54, 127, -15, -51, 127, -58, -76, 13, -10, -5, 107, 29, -112, 9, -23, -6, 2, -98, 99, -27, -107, 59, 64, 81, -60, -20, 72, 18, -93, 42, -10, -128, 127, -24, -128, 112, 113, -52, -69, -42, -17, 44, -44, 69, 8, -56, 61, -23, 70, -73, -41, 127, -22, -128, 40, 109, 27, -83, -19, -19, -72, 127, 23, -92, -75, 63, 127, 30, -128, -53, -5, -4, 127, -52, -128, 127, 71, -76, -26, -42, 42, 111, -96, -122, -12, 102, 127, 8, -128, -32, -8, -15, 55, -11, 75, -30, -107, 91, 2, -56, -2, -29, 126, 89, -88, 25, 77, -128, -6, 15, -12, 32, -90, 90, 52, -109, 34, 38, -93, 52, 127, -109, -117, 22, 74, 103, -53, 3, 0, -43, 127, -52, -42, 95, -113, -87, 89, 123, -70, -109, -40, 112, 66, -128, 9, 126, -58, 0, 127, -125, -104, 126, -38, -76, 105, 68, -128, -93, 77, 17, 49, -25, 13, 0, 37, 85, -96, -26, 24, 28, 5, -21, -12, -111, 41, 127, 7, -128, -4, 127, -110, -111, 77, 47, -7, -8, -63, 52, 37, 6, -82, -95, 127, 72, -100, 57, 7, -128, 36, 0, 72, -1, -10, 53, -110, 61, 7, -95, 77, 0, -128, 127, 30, -69, 19, 66, -89, -38, 114, -44, -32, -4, 80, -55, -78, 24, -29, 91, 17, -38, 127, -111, 4, 107, -56, -74, -14, -42, 25, 22, -72, 107, -46, 5, 26, -20, 68, -59, -22, -40, 95, 86, -52, 18, -121, -86, 11, 10, 127, 23, -128, 91, 127, -128, 17, 91, -63, -37, 20, 127, -62, -14, 55, -70, 18, -104, -42, 54, -1, 80, 6, -63, 17, 0, -77, 59, 62, -109, 107, 17, -83, 127, -89, -122, 127, 70, -37, -69, -116, 28, 44, 20, -30, 111, -51, -43, 127, -104, -128, 43, -15, 15, 127, -38, 8, 80, -128, -111, 127, 109, -100, -70, 68, 2, -11, 24, -68, -42, 114, -39, -14, -37, 21, -13, -128, 127, 122, -128, -116, 127, 36, -128, 32, -21, 52, 36, -128, 110, 104, -128, 77, 5, -60, 102, 14, -41, -56, -46, 112, 13, -75, 91, -17, -56, 41, 57, -85, -17, 100, -21, -39, -42, 36, 127, -71, -63, -15, 3, 1, 55, 42, -128, 109, -28, -51, 122, -102, 76, 64, -128, -55, -4, 100, 73, -66, -11, -53, 44, 112, 40, -128, -72, 0, 97, 17, -60, 26, 6, -62, 34, 60, -56, 102, -68, -37, 44, 19, 80, -79, -58, -61, 23, 82, 34, -61, -128, 27, 39, 97, -52, -99, 127, 15, -100, 63, 36, 55, -110, -97, -1, 82, 109, -60, -11, 81, -71, -128, 127, -25, -34, 46, -76, -17, 127, -44, -110, 127, -65, -35, 91, -77, -102, 26, 127, -23, -105, 29, 38, -56, 78, 30, -128, 41, -27, 53, 79, -92, -65, 5, 81, 44, 8, 36, -128, -39, 127, -60, -41, -27, -52, 18, 57, -7, 43, -3, 11, -72, 31, 44, -122, 110, 39, -27, -87, 59, 13, -1, -39, -45, -1, 48, -6, 12, 78, -128, 9, 37, 42, -75, -17, 127, -68, -119, 21, -22, 73, -10, -85, 104, -1, 14, 11, -105, -6, 85, 100, 0, -75, -83, -38, 80, 110, -51, -59, 1, 47, -97, 49, 83, -128, 68, 36, -38, 94, 13, -25, -32, 43, -82, -113, 52, 90, 45, -58, -75, -14, 48, 85, 54, -41, -113, -9, 70, 27, -75, -107, 81, 23, -97, 127, 35, -35, -20, 37, 86, -128, 59, 21, 11, 122, -98, -92, 66, -46, 6, 127, -68, -103, 75, -7, 12, 109, -23, -74, -8, -97, 14, 32, -106, 127, -66, -21, 97, -85, 49, -42, -39, 60, -14, 7, -38, 87, 60, -14, 72, -95, -24, 5, -1, 6, 4, 43, -72, 24, -23, -109, 90, 127, -81, -128, 97, 43, -9, -38, 6, 29, -74, -36, 58, 98, -76, 56, -14, 24, 66, -128, -21, 7, 75, -68, 24, 74, -21, -15, -85, -38, 66, 2, -119, 127, -26, -23, 37, -29, 116, 32, -128, -128, 127, 45, -48, -40, -47, -24, -8, -6, 6, 114, -1, -113, 92, 11, -32, 68, -35, 66, 22, -128, 72, 121, -128, -95, 104, 17, 56, 27, -128, 94, 65, -128, -1, 22, -11, 100, -42, -23, 82, -7, -66, -107, 113, -22, -83, 74, 46, -88, -42, 75, -55, 26, -21, -28, 76, 37, 24, -63, 68, 113, -128, -6, -10, -12, 127, -28, -70, -31, -11, 19, -66, 79, 96, -128, -86, 17, 81, 111, -113, 75, -12, -125, 96, -66, 32, 124, 2, -104, -89, 115, -26, -57, 62, -30, -34, 2, 127, 36, -30, -63, 57, 120, -128, -25, 127, -124, -9, 55, -10, 98, -108, 23, -31, -42, 127, -8, -73, -40, 78, 15, -122, -89, -34, 99, 29, -109, 99, 127, -44, -93, -54, 56, -9, -37, 28, -65, 76, -28, 0, 63, 32, 113, -113, -128, 114, -9, 45, -2, -43, 127, -128, -128, 127, -59, -56, 59, -128, 75, -2, 25, 124, -57, -109, 120, 83, -90, -99, -23, 76, 41, 32, -47, 8, -78, 2, 79, -77, 41, 78, -86, -22, 105, -56, -30, 94, -120, -3, 127, -92, 24, 17, -113, -30, 105, -37, 62, 7, -128, 36, 48, 127, -128, -128, 127, -51, 10, 127, -96, -105, 77, 9, 55, -51, -2, 55, -128, 116, 2, -22, 56, -128, 5, 95, 0, -123, 107, 51, -109, -25, 53, 127, -128, -29, 17, -15, 103, 18, 8, -128, -41, 49, 65, -30, 9, 61, -11, 48, -21, -128, 71, -1, -112, 37, 68, 70, -93, -17, 127, -22, -54, 28, -44, 46, -49, -20, 61, -128, 45, 39, -115, 127, 45, -17, -40, -93, 85, -51, -32, 30, -6, -2, 2, 64, 23, -85, -47, 123, 76, -114, -40, 27, 66, 97, -121, -123, 82, 94, -70, -100, 127, 31, -128, 44, 20, -29, 100, 60, -49, -91, -91, 127, 46, -91, 12, 77, 3, -45, 45, -103, 36, 127, -80, -49, 60, -9, 5, -52, -56, -61, 42, 44, -56, 81, 40, -4, -110, -4, 62, -1, 49, -35, -14, -86, 64, 127, -128, -72, 127, -3, 8, -22, -2, -30, -70, 64, -30, -92, 127, 58, -128, 25, 105, 3, -92, 4, 1, -6, -42, 74, -13, 12, 31, -28, -39, -85, 127, -90, 30, 62, -45, 28, 45, -54, 3, -26, -21, 127, -128, 0, 26, -55, 13, -46, -39, 79, 103, -44, -86, -86, 35, 58, 73, 65, -128, 76, -28, 0, -20, 8, 55, -63, 69, -87, -70, 41, 44, 96, -36, -35, 85, -6, -59, -85, -43, 58, 127, 53, -128, -128, 127, 37, -76, 81, -83, -8, 110, -102, -15, 91, -62, -128, 38, 127, -85, -34, 10, 3, 51, -21, 0, -46, -18, 98, 12, -68, 0, 6, -7, 12, 61, -41, -96, 29, 4, 14, 14, -69, -43, 5, -4, 56, 7, 30, 26, -31, -12, 43, -34, 44, 15, -28, -8, 3, 62, 6, -32, -126, 58, -39, -103, 93, 76, -10, -111, 127, -5, -89, 59, -80, 104, 10, -29, 127, -121, -128, 112, 24, 41, 71, -89, -88, 43, 94, -90, -72, 111, 30, -9, -59, 1, 66, 26, -113, 57, 127, -128, -90, 49, 34, -20, 114, 38, -18, 57, -80, 54, -68, -6, 85, 8, -103, 3, 47, -2, -92, -18, 103, -55, -34, 48, -60, 38, 69, -128, 127, -18, -128, 127, -11, -88, 9, -81, 127, 127, -30, -92, 37, -59, -97, 127, -80, 0, 94, -23, -8, 3, -9, -89, -41, 113, 104, -108, -1, -13, -45, 87, -63, 24, 41, -65, 121, 4, -116, 105, -11, -108, 18, -1, -3, 71, 89, -53, -88, 0, 120, 43, 0, -82, -38, 127, 19, -92, -116, 24, 52, -12, 71, -18, 43, -86, -41, 127, -79, -122, 36, 109, -83, 13, 102, -59, -73, 6, 81, -19, 0, 43, -121, 6, 114, 24, -52, -6, -65, 26, -26, -3, 6, 46, 13, -128, 127, 114, -20, -113, 36, 4, -1, -14, -128, 111, 77, -54, -73, -19, 123, 72, -20, 34, -83, -52, 61, 60, -104, 5, 80, -125, -4, 94, -79, -26, 127, -119, -54, 126, -39, -24, -47, -30, 114, -28, -112, 12, 114, -44, -8, 41, 66, -2, -111, 27, -52, -39, 56, 39, -36, -79, 115, 104, -28, 68, -85, -29, -48, 57, 51, -77, 26, 5, -72, -81, 127, -43, -70, 95, -43, -90, 127, 17, -86, 29, 12, 44, -19, -83, -99, 127, -21, 12, 48, -5, 70, -29, -42, 28, 20, 10, -15, -128, 26, 64, -30, -28, 65, -73, -116, 31, -5, 127, 4, -60, 45, -127, -9, 127, -64, -111, 127, -45, -70, -7, -41, 127, 108, -91, 29, -20, -36, -22, 43, -53, 53, 6, -76, 116, -98, -5, 100, -73, 8, -43, -89, 22, -10, 89, -23, -65, 127, 55, -76, -104, 49, 98, -128, 17, 13, 43, 127, -27, -128, -2, 127, -90, -128, 82, 127, -89, -114, 96, 71, -128, 25, 127, -128, -128, 72, 30, -22, 2, 96, 80, -111, -6, -7, -22, -38, 12, 53, -79, -4, 74, 106, -86, -6, 112, -12, 13, -128, -82, 80, 102, -49, -86, 89, 4, -43, -68, 46, 112, -75, -10, 5, 46, -66, 8, 18, -98, 20, 40, 8, -27, 112, 105, -86, -57, 66, -55, -74, 102, 6, 3, 8, -3, -55, -85, 12, 59, -8, 57, -23, -39, 36, -10, 1, -24, -3, -10, 63, -26, 25, 62, -27, -20, -19, 115, -88, -128, 70, -3, 115, 70, -128, -21, 73, -54, 41, 45, 0, 63, -96, 20, 13, -54, 3, 21, -86, 6, 7, -53, 127, 23, -128, -11, 5, 27, 63, -109, 83, 85, -81, 40, -31, -4, -26, 13, 125, 3, -97, -21, 70, -1, -7, -98, -10, 0, -104, 65, 127, -104, -128, 127, 112, -106, -109, 127, 106, -94, 48, 27, -128, 10, 30, 8, -37, 11, 55, -96, 26, 111, 65, -98, -30, 58, 0, -81, 31, 78, -22, -5, -23, 54, -70, -90, 127, -38, 35, 55, -89, 77, 46, -25, -111, -61, -10, 8, 99, 0, -55, -36, -32, 15, 23, 86, 35, 15, 30, -94, -51, 14, 54, 112, -128, 31, 11, -17, 24, -128, 44, 127, -66, -89, 112, -19, 0, 57, 21, -60, -126, 127, 44, -128, -11, 74, 102, 12, -66, -11, -75, 39, 127, -23, -42, 26, -2, -24, 6, -12, 59, -128, -65, 127, -53, -128, -12, 127, 52, 6, -115, -29, 127, -102, -2, 103, 4, -62, -34, -17, -111, 87, 15, -128, 73, 127, 66, -125, -43, 114, -128, -10, 127, -13, -17, -106, 31, 127, -128, -56, 127, -83, -87, 99, 47, -100, 23, 58, 30, -49, 9, 127, -128, -128, 127, 55, -27, 65, -28, -43, -7, -117, -47, 91, 30, 79, -20, -90, 43, 8, 37, -31, -30, -22, -116, 27, 34, 53, 85, -128, 42, 122, -128, -110, 127, -21, -48, 127, -128, -29, 92, 10, -2, 37, -55, -116, 123, 77, -24, -27, -58, 53, -58, -78, 2, -12, 98, -7, 76, -15, -93, 112, 73, -81, -3, 42, -62, -21, -15, 27, -61, -103, 48, 94, 85, -51, 8, 44, -123, 28, -19, 18, 37, -68, -62, 8, 107, -11, 37, -15, 10, -27, -87, 91, 82, -97, -45, 25, 72, -68, -126, 21, -12, 72, 75, 65, 48, -78, -39, -29, -85, 127, -55, -35, 66, -112, -28, 127, 98, -128, -19, 115, -65, 76, 11, -125, -15, 119, 85, -128, -128, 127, 27, -128, 29, 127, -49, -104, 76, 68, 11, -9, 13, -3, -13, -128, 80, 127, -128, -1, 127, -34, -81, -70, 48, 88, -49, 30, 14, 40, 76, -123, 41, -85, -31, 27, 31, 100, -86, -49, 19, -32, -53, 5, 125, 78, -128, 51, 26, -105, 43, -54, 62, 104, -128, -42, 7, 17, 127, 17, -99, 55, -60, -89, 127, 52, -68, 10, -29, 42, 107, -55, 44, -128, -4, 127, -65, -114, 27, -32, -22, 27, -75, 37, 99, -17, -48, 102, 25, -82, -25, -66, 127, 58, -128, 72, 113, -9, -115, -62, 76, -44, 82, 78, -128, 113, 11, -11, -45, 11, 127, -74, -128, 70, 127, -63, -107, -52, 45, 77, 13, -24, 42, -12, -128, 116, 10, -28, 99, -103, -56, -48, 91, -17, -3, 127, -128, 57, 109, -128, 106, 22, -26, -57, -88, 127, 38, -48, 68, -74, -116, 89, 59, 75, 30, -63, 28, -106, -47, 96, -47, 41, 45, -128, 66, 31, -17, -43, -93, 97, -32, -31, 127, -65, -85, 37, 68, -53, -5, 127, -128, 104, -14, -60, 127, -128, -75, 127, -82, -126, 74, 105, -90, -100, 127, -71, -57, 127, -112, -115, 42, 51, 35, -56, -4, 127, -25, -128, 121, -37, -34, 127, -128, -1, 116, -2, 47, -128, 56, -32, -89, 91, 43, 3, -14, 37, -28, -41, -17, 58, -14, 18, -44, -128, 127, 93, -36, -63, 4, 74, -98, 5, 31, -36, -6, -36, 9, 5, 3, 25, -55, 98, 107, -128, -43, 93, 59, -78, -128, 90, -55, 53, 69, -128, 114, -9, 9, 68, -72, 45, -45, -122, 20, 127, -12, 7, -44, -128, 18, 117, 23, -42, 62, -57, 21, -29, 46, 74, -106, -47, -56, 38, 127, -30, -57, 64, -2, -20, -54, -24, -5, 62, -1, 11, 14, 29, 8, -23, -125, 34, 88, -98, 27, -76, 81, 0, -95, 127, 43, -13, 29, 18, -128, 35, -9, 0, 56, -1, -24, 7, -32, -24, 64, -31, 18, -108, 46, -4, 26, 105, -128, -26, 11, 19, 46, 54, 13, -21, 18, -92, 4, 55, -105, 66, 46, -109, 98, -83, -61, 41, 81, 89, -128, 5, 62, -6, 86, -125, 37, 102, -18, -97, -108, 4, 79, 83, 52, -64, -82, 73, 34, -80, -92, 127, -62, -35, 56, 5, 63, -14, -111, 0, 75, -93, -34, 107, 121, -128, -128, 127, 106, 5, -128, -128, 15, 105, 124, -128, -100, 47, 103, 82, -76, 45, 49, -98, 38, -80, -44, 70, 61, 27, -122, -41, 126, 22, -127, 68, 65, -108, 36, 30, -95, 65, 32, -86, 15, -25, -17, 56, 15, -68, -47, 127, -70, 12, 66, -25, -74, 28, 37, -6, 49, -81, -15, -7, -53, 52, 20, -14, 127, 46, -128, -112, 119, 44, -10, -99, 68, -39, -36, 81, -128, 127, 15, -128, 127, 52, -8, 61, -76, -121, 99, -62, -1, 43, -97, 127, 47, -44, -45, 30, 3, 4, -89, -56, 60, 54, 31, -106, 62, -10, -58, 127, -108, 1, 7, -128, 103, -31, 76, 127, -128, 19, -40, -117, 25, 62, -29, 85, 10, -69, 108, 20, -70, 26, -42, -2, 74, -8, -77, -44, -12, 59, 56, -110, 58, 26, -30, -76, 42, 38, 59, 109, -128, 66, -19, -128, 123, -42, -65, 102, 73, 32, -36, -128, 65, 74, 37, -55, -75, -32, 56, 57, 24, -82, -8, 72, -48, -42, -35, 127, -13, -128, 98, 38, -107, 52, 78, -29, 4, 40, -91, -68, 79, 26, -25, -49, -39, 18, 52, 29, -21, -48, -58, 3, 63, -111, 88, 7, -128, 88, -36, 34, 99, 56, -85, -128, 115, 127, 0, -76, 42, -49, -128, 127, -55, 30, 38, -89, 80, -97, -10, 27, 15, 77, 28, -116, 9, 111, -128, 45, 127, -128, -77, 66, 107, -21, -92, 64, -23, -52, -5, -7, 55, 39, -109, 47, 60, -63, -42, 110, 22, -58, -58, 83, 11, -60, 127, 10, -107, -128, 100, 12, -121, 127, 73, -128, 0, -12, 51, 127, -109, 80, -80, -9, 109, -128, 36, 127, -63, -11, 52, 2, -80, 0, 80, -68, -28, 47, -45, 22, 58, 14, 27, -36, 25, -85, 25, -21, -88, 75, 69, 27, -82, 37, 11, -8, 75, -128, -11, 13, 27, 34, -128, -4, 2, 75, 73, -26, -73, 71, -14, -8, 79, 15, -12, -82, -21, -18, 57, 36, 51, -30, -85, 7, 8, -66, 9, 52, -17, -45, 76, 7, -42, 97, -45, -6, 10, -117, -27, 97, 98, -49, -69, 28, 5, -75, -80, 127, 51, -28, 24, -47, -14, -92, 123, 127, -128, -21, 6, 13, 78, 38, 53, -127, -12, 48, -128, -28, 93, -11, 65, -2, -17, -13, 31, -13, -123, 127, 83, -39, -52, -36, -80, 85, 55, -128, 43, 86, -28, 43, -57, -102, 127, -39, -28, 73, -18, 26, 34, -83, -128, 106, 66, 35, -105, -41, 22, -34, 91, -76, -24, 6, 44, 77, -99, -79, 124, 86, 0, -63, -15, -54, 30, 65, -89, 35, -47, -62, 68, -40, 14, 82, 58, -71, -64, 127, 27, -47, -38, -64, 71, 77, -63, -37, -27, 26, 62, -98, -28, 64, 32, -89, 19, 58, -20, -32, -128, 127, 48, -100, 85, 92, -128, -1, 22, -48, 105, 57, -65, -121, 37, 6, -32, -53, 127, 85, -27, -2, 24, -29, -122, 65, 73, -108, -55, 63, 12, 4, -38, 107, -68, -128, 127, -56, -128, 10, 90, 127, -127, -116, 26, 69, 40, -49, 49, -28, 79, 11, -24, 98, -13, -115, -19, 64, -30, -80, -51, -7, 76, 98, -128, 18, 127, 25, -5, -128, -108, 91, 127, -86, -65, 127, -27, 1, -43, -127, 17, 0, 81, -12, -80, 77, 24, 83, -54, -128, 8, 53, -4, 44, 127, -107, -97, 127, -37, -128, 127, 0, -45, 91, -46, -83, 71, -30, -75, 0, 4, 91, -39, 83, 66, -93, -1, -53, -3, 102, -55, 2, -42, -19, 80, -120, 73, 123, 12, -122, -128, 127, 30, -15, 20, 28, -73, -91, 8, 8, 57, -26, 94, 44, -106, 14, -41, 49, 108, -52, -6, -91, -42, 109, 38, -7, 21, -49, -29, 41, -17, -4, 9, -128, 23, -2, 59, 99, -128, 66, 97, -48, -123, 45, -1, -31, 17, -37, 49, -61, -40, 11, 8, 62, 115, -111, -90, 127, 30, -126, 1, 20, 64, -32, -100, 82, -28, -42, 127, 58, -128, 103, 10, -102, 105, 14, -103, -59, -10, 105, 27, -92, 115, 25, 1, 29, -44, -60, -13, -6, 8, -56, 24, 72, -122, 111, 106, -119, -89, 69, 127, -86, -19, -42, 45, 37, -15, -59, -55, 127, -2, 4, -94, -37, 70, -91, 3, 0, 9, 127, -46, 17, 72, 8, -112, -5, 110, -3, -93, -128, 113, 1, -52, 48, -30, -11, 93, -53, -65, 36, 70, 127, -128, -128, 124, 69, -107, 88, 61, -64, 27, 54, -21, -83, 69, 59, -95, 0, 65, -34, 21, -54, 15, -41, 1, -20, -46, 93, -106, 72, 119, -128, 42, 127, -128, -25, 37, -51, 17, 71, 66, 34, -31, -104, -9, 42, -76, 95, -1, 0, 56, 21, -22, -115, 28, -53, 25, 127, -4, -48, 45, -72, -5, 44, 51, 0, 12, -108, -7, 19, -34, 91, -128, -55, 127, 9, -57, 105, -94, -14, 94, -30, 0, 74, -115, -128, 31, 68, 123, 21, -128, -13, 127, 38, -128, 45, 78, -128, -51, 43, 30, 64, 90, -66, -128, 52, 127, -22, -76, 86, -9, -128, 98, -3, -123, 127, -11, -92, 20, 117, 108, -124, -53, 103, -83, -22, 110, -32, 13, 10, 42, -116, -69, 127, -28, -34, -4, -35, -55, 114, 6, -58, -19, -115, 127, 2, -9, 120, -62, -128, 92, 47, -82, 36, -70, 71, -34, 51, 30, -17, 94, -114, -89, 30, -3, 43, 127, -14, -128, -57, 105, 15, 34, 40, -63, -28, 83, -45, -91, 27, -1, -39, 47, 103, -52, 13, -25, -42, 55, 7, -24, -72, 93, 30, -80, 83, 102, -96, -114, 127, -12, -15, 5, -125, 30, 96, 35, -115, 60, 123, -94, -128, 89, 127, -39, -117, -35, 127, -18, 18, -59, 1, -64, 40, 24, -128, 123, 94, -51, 1, 45, -23, 11, -128, -98, 11, 124, 82, -110, 30, 21, -11, 77, -86, -19, 39, -10, -60, -13, 19, -77, 127, -24, -128, 127, -36, -47, 88, -87, -54, 54, 127, -83, -112, 30, -24, 48, 114, 49, -31, -17, -78, 0, 24, 31, -24, -114, 30, 73, 20, 6, 30, -53, 21, -72, -72, -3, 38, 127, -128, 14, 61, -128, 127, 90, -128, -54, -9, 20, -35, 119, 127, -120, -38, 26, -80, 94, 57, -55, 8, -72, -4, 4, 75, -26, -56, -2, -28, 17, -61, 74, -11, -31, 127, -80, -121, 127, 6, -128, 13, 14, -20, 127, 79, -65, -36, 37, 56, -128, 30, 28, -38, -15, 44, 30, -38, -13, -2, 121, -45, -28, -4, -12, -66, 95, 90, -128, 94, 103, -128, 64, 111, -128, 34, 41, -128, 3, 52, 52, 24, -128, 92, 127, -128, -17, 12, -14, 109, 4, -53, -83, -17, 99, 47, -90, 41, -48, -49, 92, 21, 27, -43, -11, -69, -3, 1, -68, 127, 8, 19, -25, -97, 127, -86, -31, 77, -65, -12, -34, 127, 75, -124, -37, 29, -73, 68, 27, -112, 15, 88, 93, 32, -109, -102, 127, 28, -107, -60, -4, 97, 99, -36, -128, 60, 69, -1, -91, 12, 127, -128, -1, 53, -26, -81, 56, 83, -20, -113, 14, -13, -18, 106, -11, 55, -6, -9, -60, -108, 82, 119, -128, 41, 83, -128, 61, 126, 20, -39, -19, 36, -128, -12, 61, -4, 87, -78, -62, 69, 5, -92, 63, -19, 15, 82, -128, 58, 37, -14, -55, -59, 109, -64, -57, 127, -4, -128, 127, 17, -44, 126, -128, 57, 63, -98, 82, -36, -128, 25, 3, 34, 83, 23, 46, -61, -42, -64, 2, -31, 83, 93, -93, 1, 29, 65, -36, -120, -86, 78, 56, 56, -29, -62, 104, 35, -128, 3, 8, -105, 127, -30, -38, 102, -128, 53, 7, -37, 127, -32, -37, 59, -90, -91, 63, -53, -13, 0, -10, 49, 32, 80, -93, 42, 44, -128, 89, 74, -20, 53, 1, -3, -128, 7, 62, -85, 20, 38, 99, -40, -128, 106, -15, -28, -24, 19, 106, -82, 14, 83, -5, -109, -22, 127, -109, -5, 127, -30, -89, -26, 61, -81, -57, 96, 75, -38, 46, -104, 43, 127, -128, -59, 21, 40, 53, -9, -94, -25, 99, 102, -128, -86, 127, 22, -128, -66, 24, 127, 46, -72, -25, -74, 42, 58, 15, -39, -127, 65, 47, -85, -13, 105, -2, 4, -45, 55, 127, -128, -124, 90, 127, -77, -128, 127, 127, -128, 74, 7, -128, 127, 94, -65, 52, -59, 36, 61, -128, 96, 80, -51, -128, -80, 60, 5, 70, 7, -92, 60, 48, -36, -40, 11, 77, -47, -31, 35, -8, -1, 15, -6, 82, 104, -45, -26, -106, 35, 0, -40, 126, -100, -81, 127, -30, -60, 127, 27, -25, -117, -56, 29, 3, 52, 2, 78, -6, 1, -85, 28, -10, -66, 54, -116, 86, -22, 18, 127, -31, 49, -73, -51, -48, 41, 38, -73, 11, -11, 3, -44, 31, 96, -60, 72, -51, -13, 127, -55, 19, -128, -14, 127, -49, 32, -108, -109, 11, 107, -23, -8, 127, -91, -66, 109, -56, -22, 28, -37, -36, 0, 99, -10, -98, 85, 49, -128, 103, 1, -128, 90, 31, 17, 22, 30, 39, -78, -85, 58, 22, -107, 85, -53, 40, -24, 27, 127, -58, -97, -54, 97, 82, -128, -55, -9, 93, 127, -128, 42, -45, -85, 85, -2, -74, 113, 21, -27, 28, -56, 27, 13, 62, -125, 9, 91, -128, 73, 37, -5, 117, -22, -63, 11, 62, -128, 11, 127, -25, -116, -29, 125, -21, -128, -57, 100, 116, -42, -80, -37, 97, 88, -25, -36, 3, 15, -128, 94, 40, -126, 121, -28, -105, 59, -6, -74, 88, 0, -104, 73, 37, 53, -31, 25, 94, -99, -26, 27, 54, 32, -15, -5, -27, -2, -39, -13, -18, -9, 39, -8, 89, -77, 9, -25, -11, -3, -93, 73, -36, -9, 98, 36, -128, 111, 51, -57, 4, 26, 1, -128, 104, -12, -124, 47, 127, -18, 27, -29, -128, 70, 127, -128, 2, 127, -128, -11, 120, -20, -128, -94, 127, 108, -103, 43, 18, -10, 12, -128, 26, 127, -105, -61, -23, -32, 127, 79, -20, 1, -128, 39, 27, -13, 127, -128, 3, -11, 13, 83, -60, 61, -21, -52, 20, -83, -7, 46, -83, -21, 48, 92, 104, -24, -127, -104, 127, 127, -30, -39, -2, -128, 2, 31, -128, 108, 23, 15, 89, -121, -44, 35, 99, 78, -23, -37, -128, -24, 127, -89, -47, 19, 46, 48, -36, 104, -64, -55, 100, -56, -89, 66, 13, -126, 71, 63, -27, -62, -66, 68, -24, 32, 97, -83, -32, 79, 32, 0, -128, 20, 106, -42, 39, -41, 45, 30, -126, 24, -18, -52, 127, 38, 10, -51, -42, 72, 17, -77, 15, -51, -40, 127, -28, -100, -54, -55, 127, 127, -100, 32, -12, -128, 34, -9, 13, 40, -6, 76, 15, 6, -128, -2, 86, -125, -42, 14, 110, 121, -63, -69, 109, -76, -78, 90, -18, 11, 27, -38, -9, -31, 0, -49, -12, 127, -65, -128, 36, 120, 103, -128, -13, -34, 51, 31, -128, 127, -1, -39, 115, -24, -80, 36, -56, -128, 98, 82, 42, -68, -97, 39, 57, 47, -17, -109, 43, 112, -121, 74, 75, -128, -24, 24, 0, -13, 28, 2, 127, 59, -128, 102, 37, -83, 97, -51, -10, -41, 79, 20, -104, -21, 27, 127, -17, 4, 59, -128, -31, -20, -56, 14, -24, 68, 0, -26, 47, 19, 6, -15, 81, 24, -115, -22, -53, 127, 72, -70, -55, -31, 127, -18, -58, 15, -26, -37, 25, 1, 26, -45, -46, 127, -78, -35, 30, -72, 121, 29, -20, -34, -128, 66, 127, -96, 0, 127, -119, -74, 58, 17, -112, 25, 4, 24, -3, -10, -13, -8, 127, -35, -22, -25, -64, 127, -110, -22, 53, 12, 39, -128, -9, 62, 104, -96, 9, 127, -128, -59, 25, 64, 103, -89, -102, 115, 114, -111, -92, 127, -92, -97, 115, 38, 60, -128, -8, 127, 13, -128, 15, 55, -110, 0, -61, 3, 56, 127, -99, -51, 65, -72, 49, -51, 35, 127, -128, 8, 18, -28, 109, -105, 95, 23, -128, 127, 36, -32, 109, -94, -128, 93, 119, -62, -128, 69, 121, -87, 8, 65, -128, 80, -12, -91, 22, 28, 28, -104, 36, 15, 54, 96, -57, -8, -66, -31, 105, -23, -28, -7, 77, 10, -106, 17, 127, -63, -107, 77, 80, -105, -78, 127, -71, -80, 72, -41, -54, 69, 42, -66, 117, -65, -116, 65, 83, -37, 31, -7, -17, -6, -8, 57, -30, 108, -125, -32, 45, -39, 42, -91, 52, 127, -128, 29, 55, -77, -18, 6, -8, -7, 127, 58, -41, -128, -20, 44, 8, -31, 47, -14, -31, 32, 44, -27, -79, 120, 80, -40, -74, -61, 60, 127, -128, -45, 127, -91, -87, -59, 116, 44, -73, 87, -41, -108, 95, 82, -64, -89, 57, 127, -114, -128, 11, 126, -14, -74, 88, -80, -109, 127, 2, -49, 127, -105, -64, 95, 4, -9, 34, -75, 75, -10, -128, 43, 39, 72, 86, -30, 10, -19, -13, -97, 9, 127, 22, -128, -77, 117, -90, 1, 55, -42, -17, -28, 53, 63, 22, 90, -108, -92, 58, -65, 60, 37, -66, 127, -52, -128, 127, -76, 49, 85, -128, 92, 44, -128, 87, 116, -60, 27, -43, -128, -8, 97, -34, 42, -35, 32, 122, -128, -21, -40, -7, 127, -47, -39, 114, -60, -128, 34, 96, -95, -97, 127, 127, -58, -128, 78, 59, -27, 66, -15, 42, -128, -60, 14, 55, 87, -128, -1, 127, -23, -48, -21, -27, 127, -71, -92, 77, -18, -60, -42, 87, -17, 83, 28, -36, -52, -75, 29, 111, -14, -128, 127, 1, -79, 127, -99, -128, 30, 94, -41, 17, 39, -60, 24, -49, 69, 78, -11, 48, 6, -27, -26, -128, 62, 127, -45, 3, -72, -128, 121, 66, -128, 54, 75, 2, -6, -13, 43, 18, -116, 46, 24, -71, -14, 18, 61, 43, -61, -99, 127, -53, -115, 74, -11, -56, 17, 127, 94, -99, 17, 13, 6, -93, -114, 93, 63, 61, -117, -32, 82, -37, -26, 79, 74, -52, -59, -8, -2, 31, 79, -105, 27, -46, -23, 9, -96, -11, 127, -8, -106, 127, 10, -100, 44, 80, -17, -49, -6, -95, -77, 47, 25, 79, -68, -40, 32, 29, 96, 24, -96, 25, -35, -98, 127, 86, -91, -128, 117, 57, -128, 46, 6, 48, 126, -128, -15, 127, -128, -12, 25, -108, 127, 6, 7, -83, 9, 31, -52, 127, -128, -99, 127, -8, -14, 75, -64, -104, 121, 7, -35, -40, 19, 127, -128, 4, 49, -12, 109, -128, -27, 98, -18, -43, -35, -6, 68, -70, 29, 51, -128, 99, 93, -28, -69, -68, 54, 20, 15, -59, 77, -29, -98, 127, -62, -52, 89, -5, -28, -23, 57, 122, -121, -102, 85, 1, 40, 108, -36, -87, -26, 44, -36, 76, 8, -98, 6, 30, 109, -25, 6, -13, -13, -59, -102, 122, 28, -13, -76, 6, 127, -24, -62, 26, 52, 10, -128, -51, 122, 25, -128, -85, 76, 13, -48, 58, 99, -53, -69, 58, -37, -54, 17, 109, 30, -86, 35, 106, -111, -34, 106, 30, -27, -128, 102, 25, -122, -55, 127, 127, -74, 23, -98, -128, 43, 10, 64, 103, -46, 27, -37, -41, -37, -13, 65, -40, 121, -99, -76, 10, 57, 22, -128, 39, 37, 114, 24, -91, 86, 0, -91, 56, -8, -26, 63, -8, 14, -32, -56, 11, -40, 107, -74, -66, 87, -6, -72, -12, 94, -7, -4, -40, 22, 40, -48, 91, -6, -128, 43, 47, -15, 127, -91, -128, 115, 127, 6, -64, -47, -42, 102, 95, -128, -113, 32, 112, 25, -44, -60, -24, -46, 93, 80, -30, -23, -114, 66, 124, -106, -80, -10, 111, 10, -128, 127, 78, 28, -23, -128, -15, 126, -36, -100, 3, 6, 78, 110, -125, -112, 56, 7, -8, 109, 81, -6, -114, 10, 53, -22, 94, -75, 1, 5, -24, -99, -48, 103, -103, 89, 115, -121, 22, 85, -41, 17, -66, -109, 127, -32, -71, 127, -30, -53, 95, -98, -19, -17, -77, 2, 127, -27, -63, 127, -14, -95, 63, -71, 9, -6, -128, 127, 25, 42, 23, -128, 65, 112, -79, -30, 85, 65, -82, -92, 57, -22, 8, -1, -66, 115, -6, -102, 127, -42, -128, 119, 59, -110, 57, 62, -115, -71, -22, 110, 115, -42, -14, 18, -80, -55, -10, 13, -15, 69, 68, 35, -112, -68, 34, 15, 2, 35, -48, -91, 127, 0, -128, 64, 120, -117, -51, 14, -29, 71, 120, -72, -116, 109, 99, -13, -128, -52, 6, 0, 127, 69, -123, -95, 6, 69, 66, 6, -87, 18, 127, -97, -122, -25, 125, 127, -128, -119, 127, 3, -53, 92, -65, 47, 1, -107, 39, 18, -9, 1, 49, -9, -74, -68, 52, 77, -3, -34, -104, 127, -25, -128, 51, 5, 7, -14, -29, 59, 11, 94, 57, -12, 24, -128, 79, -9, -65, 74, 14, -43, -107, 75, 105, -36, 1, 0, -105, 4, 120, -20, -87, 103, 12, -79, 107, 10, -63, -119, 76, 127, -34, -24, -31, -7, 12, 2, -11, -21, -106, 12, 92, -68, 87, 1, -59, 82, -35, 56, -112, -56, 38, -3, 6, 20, 127, -87, -110, 75, -13, -40, 23, -38, 93, 127, -54, -52, -3, -59, 83, 34, -47, -19, 10, 28, -14, -17, -75, -1, 7, -26, 91, 2, 0, -65, -122, 127, 1, -44, -8, -2, 98, -32, -9, 28, -44, -19, -54, 109, 105, -128, 2, 58, 5, 7, -96, 38, -40, -9, 127, -76, -1, 77, -29, -10, 14, -121, -48, 25, -7, 89, 18, -68, -90, 13, 120, 14, -48, 95, -37, -94, -26, -66, 126, 125, -64, -124, -19, 86, 44, -27, -128, 88, 13, 29, 71, -128, -42, -8, 34, 95, 78, -128, 32, 127, -128, -5, 32, -128, 59, 127, -85, -10, 122, -122, -30, 59, -54, -56, -32, 0, 74, -19, 43, 120, -128, -68, 127, -47, -79, -1, 92, -11, -128, 127, -71, -35, 112, -70, 44, -29, -57, 0, -34, 37, 40, 83, 53, 18, -128, -125, 25, 96, 1, 68, 20, -106, 29, -39, 46, 91, -43, -53, 80, 39, -128, 58, -6, -14, 20, -128, -32, 121, 3, -108, 127, 72, -128, 59, 96, -128, 85, 76, -35, -76, -1, -7, -23, 127, -54, -128, 82, 94, -4, -32, -11, -89, -9, 127, -128, 21, 29, -128, 127, -2, -58, 57, 74, -27, -77, -11, 41, -41, 75, 0, -111, 71, -44, 91, 12, -89, 127, 83, -128, -9, 58, -9, 83, -128, -7, 127, 22, -22, -9, -38, 19, -79, 25, 88, -102, -54, 43, 123, -100, -72, 127, -28, -48, 120, -128, 7, 20, 7, 85, -128, 28, -43, -91, 80, -28, 85, 14, -128, 69, 127, -2, -108, -61, 29, 127, -18, -29, 24, -44, -91, -42, 57, 38, 96, -56, -51, 93, -34, -7, -45, 74, -27, -79, -19, 21, 79, 21, 30, -40, -72, 44, -36, -22, 127, -12, -42, -38, 0, -49, 79, 55, -98, -21, -51, 4, 75, 80, -98, -100, 76, 52, -66, 21, 127, -96, -114, 86, -35, -76, 17, 55, 113, -25, -126, 97, -36, 27, 14, -28, 8, -88, 37, 69, 39, -58, 105, -47, -123, 13, 8, 102, 20, -25, -34, -6, 74, -3, 38, 32, -52, -105, -57, 66, 22, 3, -69, 35, 20, -47, 4, -1, 51, -2, 65, 79, -34, 12, -128, 39, 127, -128, -11, 4, 20, 95, -8, -63, -58, 71, -24, -128, 127, 62, -78, -2, -116, 48, 127, -128, 36, -18, -96, 76, -18, 0, -30, -3, -22, 15, -4, 117, 49, -26, -36, -78, 112, -80, 53, 47, -128, 35, 100, -66, -80, 32, 89, -52, 80, 71, -128, 110, 15, -18, -49, 46, -28, -75, 40, -82, 125, 24, -123, 29, 4, -1, 100, 71, -49, -3, -69, -3, -12, 3, 117, -128, 72, 5, -128, 127, 40, -72, 18, 106, -100, -25, 127, -123, -104, 127, -21, 14, -14, -100, 39, -43, 86, 92, 59, -126, -57, -2, 28, 75, -1, -49, -22, 64, -79, 52, -22, -27, 127, -14, -79, -91, 3, 35, -51, 49, 127, -42, -92, -53, 53, 89, -103, -20, 35, -36, 10, 124, -45, -113, 13, 127, -22, -9, 18, -57, 31, -2, -54, 8, -5, 23, 66, -42, 53, 42, -128, 53, 6, -87, 127, 14, 32, -114, -128, 74, 3, 48, -31, -30, 114, -23, -78, 127, -42, -54, 71, -4, -62, 23, -2, -62, 45, 28, 116, -97, -107, 127, 97, -106, -88, 98, -46, -87, 127, -51, -13, -41, 3, 127, -83, -36, -77, 72, 51, -110, 15, 90, 68, -52, -77, 71, 63, -42, -53, -3, 52, 19, -41, 8, -83, 66, 61, -125, 17, -15, 60, -45, -47, 62, 56, 56, -23, 9, -28, -128, 95, 127, -71, 5, -74, -105, 45, 127, -2, -12, -9, -100, 46, -44, -124, 127, -20, -51, 35, -36, 121, 47, -49, -89, -39, 44, -29, -52, 27, 98, -24, -69, 46, 99, 82, -71, 25, -34, -69, 63, -45, -68, -63, 127, 32, -128, 127, 19, -57, 120, 13, -98, 21, -29, -29, 127, -24, -62, 70, 35, -128, 52, 127, -124, -5, 78, -128, 25, 11, -24, 49, -60, 91, -19, -89, 126, 7, -128, -34, 127, 109, -25, -110, -14, -53, 55, 73, -71, 24, -39, -30, 56, 5, -68, -24, 6, -17, -18, 127, -48, -6, 30, -64, 74, 13, -124, 15, 31, -122, 127, -17, -128, 127, 30, -23, 86, -71, -95, 20, 111, 9, -14, 9, -128, -77, 127, 21, -102, -27, 15, 83, -83, 58, 10, -3, 66, -106, 10, 62, -2, -56, 51, 60, -111, -63, 82, -56, 27, 127, -42, -18, -7, -13, -40, 21, 91, -93, -98, -4, 37, 66, 34, -9, -73, 90, -24, 0, -22, -6, 59, -60, 127, -89, -128, 53, 4, 92, -47, 69, 23, -46, 39, 21, -66, 1, 74, -128, -79, 127, -18, -45, 9, 22, 124, -70, -79, 106, 108, -112, -55, -19, 62, 58, -128, 110, 62, -95, 1, 58, -36, 26, 43, -128, 59, 127, 8, -95, -19, 112, -8, -5, -96, -128, 22, 127, -69, -62, 127, -128, 59, 32, -128, 121, 56, -72, 34, -64, 66, -12, 0, 60, -128, 55, 34, 73, -10, -103, 18, -26, 14, 19, -60, 82, 19, -39, 72, -8, -71, -14, 80, -55, -8, 107, 53, -110, -110, 89, 21, -88, 87, 14, -21, -89, 72, 44, -128, 71, 100, -34, 41, -76, -7, 127, -3, -128, -25, 74, 2, 49, 52, -75, -128, 83, 38, -128, 127, 73, -41, -40, 28, 35, -18, 1, -47, 52, 9, -24, -73, -69, 127, 110, -128, -28, 125, -128, 19, 55, -72, 53, -78, -9, 127, -83, 32, 127, -128, 10, 52, 1, -38, -97, 47, 100, 48, -5, -5, -86, -23, 75, 28, -82, 40, -82, -107, 127, -35, -127, 127, 79, -119, 76, 97, -128, -128, 127, -12, -128, 127, 51, -128, 71, 127, -106, 13, 36, -72, 9, -42, -85, 57, 127, 19, -128, 72, 92, -4, -128, 8, 127, -77, -76, 39, 28, -68, 71, -28, -37, -39, -109, 127, -41, -40, 127, -107, 4, -34, 59, -29, -105, 127, 17, -115, -8, 115, -53, -96, 117, -20, -89, 46, 97, 12, -109, -18, -9, -70, 114, 103, -128, 41, 115, -128, 32, 43, -23, -10, 19, 30, -38, -53, 4, -13, 23, -6, -116, 127, 75, -128, -31, 127, 34, -128, 51, -69, 7, 127, -128, -30, 100, -69, 3, -5, 12, -11, 48, -15, -20, 99, -128, -10, 14, -5, 124, -1, -19, 35, 2, -92, -116, -23, 58, 76, 32, -125, 56, 34, 25, 127, -128, -15, 64, -1, -26, -105, 35, -13, 78, -26, 57, 89, -47, -86, -62, 78, 104, -88, -64, 119, -22, -30, 49, 66, -113, -100, 127, 83, -72, 9, 27, -39, -14, -87, -29, 114, -41, -34, 97, 26, -32, -6, -29, -74, 65, 52, 1, -26, 4, -36, -92, -7, 86, 127, -128, 21, 34, -28, 98, -35, 11, -60, -25, -35, 14, 94, 35, 4, -104, -15, 71, -128, -12, 8, -8, 7, 73, -13, -11, 75, -81, 80, 56, -128, 38, 112, -128, -106, 90, 127, -128, -76, 102, -19, 72, -78, -70, 127, -110, 26, 91, -31, -72, -128, 127, 60, -128, 55, 87, -121, -57, 49, -34, -31, 99, -35, 54, 127, -128, -9, 110, -70, -92, -5, 111, 121, -91, -113, 85, 29, -96, -3, 7, -13, 41, -43, 56, 83, 5, -53, 6, -58, -35, 127, -95, -128, 127, -13, -128, 19, 127, 85, -57, -117, -70, 98, -28, 1, 127, 49, -126, -111, 53, 40, 23, 49, 27, -82, -10, 36, 60, -47, -15, 60, -112, 83, 108, -128, -109, 127, 15, 21, 26, -34, 83, -52, -93, -94, -5, 5, 117, 12, -107, -21, 60, 95, 23, -107, 56, 1, -63, 111, -44, -43, -55, 81, -3, 24, 121, -124, 1, -12, -62, 30, -40, 31, -48, 27, 87, -98, 69, 8, -78, 127, -59, 17, 39, 3, -61, -87, 10, 70, -21, -22, 19, -70, 52, 17, -7, -47, 93, 127, -66, -123, -18, 88, 49, -69, -75, 127, 10, -11, -43, -22, 122, -103, 26, -21, -89, 123, 36, -80, -2, 59, -109, -14, 127, -66, -128, -18, 75, 125, -114, 19, 127, -128, -45, 47, -20, 57, -4, -128, 52, 105, 9, -22, -128, 43, 109, -43, -28, 0, -83, -25, 32, -34, 127, -27, -53, -14, -39, 20, 73, 66, -128, 75, 115, -23, -73, -45, 40, 76, -11, -104, 39, 4, 26, 85, -128, -3, 43, 19, -46, -29, -7, -49, 127, -99, -28, 98, -109, -70, 87, 127, -51, -38, 64, -83, -18, -43, 65, 14, -128, 63, 70, 38, 62, -60, -26, -44, -62, 26, -52, 52, 127, -66, -128, 122, 25, 3, -10, -72, 112, 65, -78, -88, 71, -48, 26, 8, -81, 91, -9, -6, -44, -87, 76, -18, 52, 5, -52, -12, 1, 79, 32, -45, 14, 98, -125, -100, 109, 18, 9, 25, -61, -27, -56, -22, 124, -73, -1, 36, 19, 18, -128, -13, 89, 68, -35, -48, 80, 92, -72, -76, 25, -36, 69, 34, -117, -48, 127, -52, -20, 127, -24, -46, -114, 119, 73, 3, -112, -74, 45, 65, 89, -114, -103, -4, 127, 3, -60, 71, -53, -88, -36, 127, 59, -128, -13, 127, -25, -114, 92, 127, 9, -91, -62, -64, 34, -17, 100, 68, -98, -10, -10, -2, 31, 30, -9, -12, 75, -42, -126, 31, 23, 25, -68, 92, 45, -88, 35, 22, 13, -73, 13, 29, -4, 97, -36, -128, 124, 53, -91, 23, 9, 80, 9, -114, -34, 1, 68, 0, -69, 127, -15, -9, -43, -39, 72, 3, -95, -75, 36, 76, -3, 44, -49, -128, 127, 66, -128, 42, 127, -6, -128, -3, 79, 32, 26, 38, -124, -49, 41, 3, 36, 35, -11, -5, 27, -124, 7, 90, -54, 41, -28, -12, 81, -115, 58, -8, -4, -46, -128, 127, 98, -99, -65, 32, -26, -31, 44, 11, 63, 79, -128, -45, 117, 36, -54, -71, 110, 127, -128, -86, 127, -12, -105, 73, -85, -40, 38, 74, 57, -117, 53, -26, -21, 127, -38, -12, -98, 49, -10, -28, 124, -128, -39, 20, 85, 46, -56, 40, -8, -2, -56, -11, -9, 34, 18, -85, -12, 62, -11, 12, 127, 30, -128, -39, 127, -13, -96, 77, 30, -106, 83, -71, -19, -4, -39, 59, 43, -64, -85, 45, 90, 8, -9, 111, -119, -128, 32, 26, 70, 14, -119, 53, 48, -98, 10, -2, 83, 94, -122, -26, -4, 120, 46, -30, -42, -128, 34, 127, -57, -51, 8, 72, -14, -128, 127, 19, -128, -1, 57, 119, -34, -25, -25, 21, 59, -62, 49, -13, -128, 124, 99, -128, 87, -3, -128, 11, 20, 36, 127, -42, 11, -18, -128, 127, -24, -128, 28, 35, -9, 85, -42, 0, 48, -61, 18, 73, 97, -128, -88, -8, -38, 127, 12, -128, -11, 60, 13, -36, 127, -55, -35, 127, -72, -128, 100, 103, -128, 90, 127, -128, -25, 127, -110, -128, 78, 61, 100, -57, -22, 6, -103, 127, -60, -41, 9, -66, 17, -7, 83, 100, -30, -108, 51, 88, -81, -40, 7, -9, 43, -80, 86, 7, -128, -13, 5, 93, 45, -89, 80, 12, -80, 12, -42, 58, 117, -76, 26, -66, -39, 100, 40, -78, -5, 124, -128, -38, 52, -7, 100, 52, -56, 28, -124, 8, 127, -124, -51, 13, 20, -19, 38, -61, -38, 127, -13, -79, -41, 14, 45, -89, -63, 93, 24, -72, 0, 47, 35, 8, 71, -26, -88, 58, -32, -13, 64, -98, 99, -35, -73, 115, -48, -41, 55, -56, -44, 51, 22, 57, 63, -123, -24, 127, -39, -128, -75, 127, 35, -46, 7, -39, -68, 78, 127, -108, -90, 41, 26, -38, 17, -47, 44, 127, -95, -91, 102, 38, -49, -34, -48, 15, 34, -80, 17, 4, -76, 92, 116, -9, -112, -58, 127, -38, 17, 114, -106, -40, -64, 122, 61, -55, -83, -38, 102, -25, 54, 7, -128, 10, 127, -32, 25, -29, -70, 37, -56, 37, 120, -98, -119, 9, 38, -15, -18, 53, 66, 63, -35, 31, 23, -119, -15, 93, 26, -110, -74, 87, 51, -19, -97, 37, -8, -103, 127, 66, -71, -45, -41, 54, 13, -9, 23, 45, 0, -128, -44, 73, 61, 103, -90, -60, 23, -105, 43, 23, -53, 115, 105, -128, -48, 12, 35, 87, -96, 51, -27, 27, 127, -76, -76, 11, -45, -45, 31, 116, -56, -14, -5, 48, 76, -91, -12, 70, -11, 24, -103, -20, 127, -34, 45, -128, 26, 70, -63, -32, -103, 127, -14, -128, 75, 66, 26, -10, 14, 89, -95, 3, 63, -99, 83, -46, -128, 77, -8, 41, 56, -106, 52, 2, -90, 61, 43, -69, -47, -9, 56, 0, 90, 32, -104, -29, 107, 100, -52, -35, 40, -107, -25, 72, -6, 18, -6, 68, -105, -128, 115, 106, -73, -62, 119, 13, -6, -28, -48, 125, -49, -128, -21, 46, 41, 19, 10, -9, -29, -1, -38, -15, 53, 80, 49, -111, -45, 49, 114, -4, -112, 75, -88, 43, 3, -128, 68, 127, 6, -128, 95, 127, -128, -119, 14, 94, 45, -13, 81, 5, 15, -128, 32, 58, -69, 77, -52, -83, -55, 73, 64, 19, -85, 25, 56, -113, 61, 114, -116, -116, 127, 124, -7, -11, 32, -128, -62, 80, 22, 12, -93, 44, 51, -103, 113, -23, -19, 59, -128, 113, 85, -39, -68, 44, -23, -8, -37, -128, 116, 0, -74, 24, 127, 127, -128, -14, 127, -66, -127, 14, 127, -40, -128, 5, 90, -65, -6, 68, -41, 75, -19, -98, 37, 109, -98, 24, 97, -128, 65, 127, -128, 19, 31, -128, 127, 3, -15, 98, -18, -116, -70, 127, 0, -52, 96, 85, -90, -70, -34, 102, -43, -42, -2, 0, 59, -95, 23, 123, -40, -106, 108, 20, -128, 109, 53, -128, -28, 42, 86, 98, -80, -128, 44, 112, -9, -55, 55, -98, 66, 14, -128, 34, 127, -32, 31, -5, -88, 87, -105, 71, 123, -2, -66, -128, 112, 127, -128, -107, 3, 127, 127, -82, -128, 30, 35, -7, 125, 47, -74, 34, -125, -15, 24, -25, 127, -128, 15, 81, -128, 127, -46, -128, 127, 40, -120, 57, 1, -64, 91, 0, -77, 39, 108, -53, -121, -40, 127, -5, -128, 127, -7, -102, 87, -14, 97, 25, -128, 108, 72, -52, 7, 30, 15, -55, -73, -58, -29, 90, 27, 20, 82, -22, -97, 6, 120, -77, -35, 97, -81, 9, 5, -78, 92, 45, -61, 30, -116, 24, 91, -38, 3, -89, 41, -10, 17, 117, -114, 23, 7, -46, 72, -93, -59, 127, 97, -128, -95, 107, -73, 23, 71, -60, -22, -20, -9, 111, -31, -115, 127, 60, -119, -88, 127, 64, -107, 36, -4, 12, 10, 8, -1, -99, -78, 127, 22, -128, 6, 85, 91, -73, -45, -20, 62, 76, -85, 89, -12, -76, 1, -68, -4, 37, 30, -61, 113, 103, -35, -49, -32, 15, -35, -62, 74, 74, -128, 107, 94, -128, 38, 2, -39, 127, -23, -128, 22, 126, -90, 20, 46, -121, 127, -5, -46, -29, -22, 55, 79, -63, 10, 39, -41, -29, -14, 29, 7, 44, -58, -77, 76, 121, -80, -117, 71, 87, -69, -98, 34, 36, 68, 37, -52, 44, -114, -93, 127, 8, -40, 55, -14, -2, -88, -45, 126, 40, -22, -23, -59, -79, 91, 10, -128, 20, 52, 82, 64, 14, -128, -46, 53, 81, -15, -128, 127, 24, -83, 75, 78, -97, -53, 73, 55, 42, -128, 39, 86, 0, 8, -128, -29, 69, 15, -17, 44, 99, -96, -36, 116, -81, -90, -9, 9, 52, -37, 107, 70, -94, 24, -35, 4, 112, 31, -93, -32, 92, -64, -126, 103, 103, -128, 70, -24, -78, 42, 26, 14, -52, 25, -90, 66, 81, -128, 75, 125, -128, 23, 6, -10, 0, -17, -11, 119, 7, -105, 121, -121, 30, 127, -23, -22, -128, 53, 110, -81, 92, -58, -22, 34, -68, 109, -95, -128, 127, 125, -85, 49, -52, -32, 27, -45, -56, 22, 65, -45, -45, -34, 32, 127, 95, -128, -79, 127, 87, -128, -85, 127, -30, -109, -4, 127, -45, -128, 127, -80, -128, 117, 123, -17, -111, 10, -60, 27, -7, -21, 127, -102, -24, 39, -120, 76, 48, -14, 22, -43, 11, 121, -95, 29, 0, -94, 127, -42, -128, 127, 72, -128, 63, 15, 20, 97, -18, -4, -74, 14, 1, -93, -38, -55, 109, -7, -19, 127, 4, -128, -36, 22, 116, 52, -128, -28, 1, -12, 86, 0, -106, 127, 19, -53, 25, -110, 85, 9, -109, 20, -1, 54, 77, -83, 34, -12, -52, 42, -44, -37, 42, 64, -15, -32, 123, 19, -70, -71, 49, 9, -107, 127, -59, -39, 110, -69, 76, -42, -9, -43, -15, -18, 18, 55, -96, 51, 8, 39, 49, -41, 29, -70, -122, 15, 92, -42, 44, 15, -108, 93, -8, 9, 23, -23, 2, -92, 127, 29, -125, 127, -6, -128, 116, 4, -87, 18, 23, 107, 46, -85, -80, 83, 3, -56, 97, -100, -55, 127, -120, 61, -9, -79, 65, -18, 83, 19, -74, 28, 89, -128, -26, 89, -123, 49, 65, -25, 57, -68, -64, 110, 1, 38, -2, -128, 25, 58, -43, -31, -26, 75, -18, -25, -10, 48, -11, -111, 75, 105, -85, -53, 127, 34, -8, 42, -79, -92, 61, -54, 1, 127, 48, -128, 35, 48, -103, 58, -109, 53, 127, -128, -25, -32, 27, 108, -23, 8, 23, -107, -69, 127, 19, -128, 19, 55, -119, 103, 108, -63, -111, -34, 86, 92, -5, -75, -4, -64, -51, 82, -13, -99, 127, 100, -128, 13, 20, 66, 13, -128, -32, 127, -46, -2, 3, -21, 46, -113, 116, -65, 22, 127, -107, -48, 89, -73, -117, 57, 24, -19, 100, 3, -88, 44, 107, -9, -128, -12, 63, 30, -1, 28, -23, -4, 15, -14, -27, 27, 97, -128, 9, 111, -2, -65, -122, 97, 19, -90, 114, 37, -78, 18, 43, 51, -128, 9, 42, -81, -47, 117, -56, -42, 127, -78, -14, -27, -88, 127, -6, -128, 7, 127, 126, -128, -49, 9, 64, 114, -86, 21, 2, -125, 41, 57, -105, 105, 22, -51, 17, -19, 59, -37, -25, -22, 83, 105, -94, 31, 56, -94, 42, 53, -92, -13, 59, 0, -9, -34, -36, -52, -44, 127, -29, -5, -9, -91, 93, -19, 44, 61, -5, -58, -121, -25, 77, 112, 34, 14, -17, -58, -40, 27, 1, -126, 23, 29, 73, -30, 6, 30, -80, -2, -61, 89, 127, -76, -128, 43, 95, 69, -91, -52, 15, -53, 66, 88, -99, -44, 105, 75, -109, -114, 113, 46, -52, -97, 125, 10, -122, 127, 9, -14, 79, -19, -85, 29, 95, -60, -123, 48, 9, -17, -42, 0, 112, 18, -108, 56, -36, 3, 125, -128, -74, 15, 104, 13, -83, 38, 26, 15, -71, 86, -8, 14, 59, -91, 76, -27, -128, 111, 127, -128, -59, -62, 95, 3, -34, -14, 27, 112, -18, -39, -23, 87, -32, -73, -82, 79, 106, -58, -102, 80, 17, -104, 88, 78, -128, -18, 57, -114, 91, 3, -12, -17, -47, 80, -45, 100, 54, -128, 68, 39, -24, 38, -54, -47, 120, 46, -128, 83, -8, -71, 124, -23, 46, 11, -90, -72, -37, 127, -37, 12, 127, -60, 22, -78, -128, 20, -8, 86, -5, 19, 120, -3, -104, -83, -7, -15, 125, -23, 28, 110, -66, -9, -62, 24, -28, 8, 97, -73, -18, -89, -14, 77, 49, -31, -27, 107, -60, 0, -6, -26, 46, -70, -20, 102, -8, -34, -68, -72, 127, -49, -128, 116, 94, -21, -55, -80, 31, 10, 9, 127, -83, -128, 53, 127, -11, -128, 85, 120, 11, -117, -47, 60, 3, -75, -18, 5, 48, 59, -69, 27, 10, 7, -55, -36, -7, 48, 32, -15, 53, 75, -53, -24, 94, -9, -21, -105, 52, 53, -128, 74, 89, -28, -56, -85, 91, 66, -81, -52, 127, 27, -32, -9, -128, 107, 94, -128, -36, 127, 5, 9, 13, -7, 11, -78, 29, -44, 15, 41, -23, 73, -83, -75, 49, 12, 22, -49, -99, 127, 77, -128, 19, 48, -19, 56, -35, -105, 94, 70, 23, -58, -69, 77, -64, -51, 8, -62, 65, 127, -26, -112, 61, 80, -7, -83, -46, 20, 19, 37, -38, -87, 107, -66, -26, 80, -5, -68, -15, 81, 7, 1, 24, -29, -105, -28, 77, 48, -98, -9, 37, 66, 57, -98, 6, 51, 9, -45, -111, 77, -44, 46, -11, -128, 127, 103, -79, 14, -114, -51, 60, 89, -57, -93, 70, -8, 65, -82, 51, 127, -103, -70, 69, -44, 24, 70, -128, 82, -12, -87, 115, -47, -43, 68, 19, -64, 25, -14, -81, 73, 78, -22, -28, 26, 68, -7, 54, -65, -49, 127, -106, -108, 69, -69, 47, 54, -30, 96, -100, 4, 2, -15, 127, -51, -103, -22, 80, 69, -82, 34, -57, 39, 1, -80, 60, 71, -56, -72, 48, -99, 31, 106, -57, 61, 28, 17, -45, -128, 120, 9, 3, 117, -128, -1, 68, -76, -29, -29, 2, 45, 127, -61, -68, -31, 48, 127, -128, -128, 105, 49, -97, 97, 127, -128, -2, 27, -65, -85, 81, 9, -69, 121, -98, 3, 76, -57, 114, -2, -56, -44, -102, 99, 51, -23, 59, -53, -35, 98, -59, 66, -47, -117, 127, -125, -7, 127, -86, -80, 66, -9, -64, -4, 80, 20, -7, -39, 6, 96, -35, -51, 14, 83, -128, -74, 66, 64, 17, 29, -31, 1, 87, -77, -80, 57, 30, -98, 23, -47, 15, 49, -83, 127, 34, -128, 9, 27, -5, -26, 127, -47, -72, 127, 0, -4, -127, -74, 66, 48, 100, 27, -108, 41, -46, 7, 55, -9, -55, -128, 127, 103, -99, -95, 55, 127, -78, -126, -23, 106, 29, -119, 69, 127, 18, -85, -51, 88, -18, 9, -21, -63, 40, 65, -65, 2, 68, -4, -13, 14, -115, -54, 127, -61, 32, -6, -113, 127, 7, -128, 63, 40, -40, -66, 35, -14, 6, 127, 28, 19, -18, -128, -3, 26, -107, 127, -13, -28, 120, -20, -20, 5, -42, -75, -44, 127, 62, -128, 107, 72, -80, -24, -65, 75, 54, -75, 91, -103, -90, 127, -76, -128, 127, 70, -128, 110, 0, -124, 71, 122, -112, -128, 127, 3, -62, 90, -40, 2, 127, -128, -64, 73, -3, 51, -47, -95, 21, 12, -36, 79, 127, -119, -25, 119, -46, 41, -9, -2, -54, -123, 127, -11, -68, 36, -2, 91, -112, 4, 88, 0, 93, -128, -68, 94, 31, 29, -3, -128, 49, 127, -65, -12, 62, -63, -82, 59, -20, -81, 28, 83, -17, -72, 82, 94, -46, -74, -3, 70, -78, -99, 119, -22, -77, 6, 82, -51, 43, 73, -128, 127, -11, -19, 104, -128, -35, -9, 88, 90, -97, -36, -7, 76, 70, -121, 28, 24, -2, 20, -83, -76, 116, -8, -88, 32, 3, -10, -11, 45, 25, 24, -64, 62, -1, 7, 113, -46, -128, 56, 46, -62, -25, 48, 11, 8, 127, -128, -108, 127, 18, -46, 75, -59, -11, -22, -20, -9, -65, 127, -12, -3, -20, -34, 47, -18, 4, -22, -58, 40, -6, -39, 127, -42, -128, 28, -28, 127, 14, -128, 121, 36, 31, -3, -128, 26, 127, -40, 10, -92, -30, 3, 60, 94, -36, -47, -70, -24, 88, 20, -24, 74, 12, -58, 37, 46, -79, 44, 6, -23, -66, -59, 57, -27, -91, 54, 127, 32, -128, -27, 127, -29, -30, 40, -86, -22, -39, 6, 102, 2, 58, -85, -68, 73, 47, -36, -63, 13, 10, -45, -37, 106, 39, 17, -119, -7, 61, 31, 20, -76, 35, -30, -61, 9, -18, 14, 127, -64, -128, 53, 127, 66, -38, -91, -5, 11, 63, -74, -128, 85, 32, -4, -42, 122, 2, -128, 108, 66, -91, -55, 0, 103, 59, -63, -79, 47, 127, 9, -21, 28, -99, -36, 127, -128, -117, 99, 76, -92, -2, 110, -56, 65, -95, -54, 127, -128, 15, 51, -12, -80, -36, 127, 10, -128, -77, 124, 97, -128, -10, 115, -108, -105, 89, 2, -78, 122, 61, -8, 56, -105, -48, 44, -74, 51, -11, -114, 127, -42, -53, 127, -122, -54, 91, 89, -42, 7, 55, -94, -91, 48, -5, -36, 94, 42, -40, 42, 2, -128, 77, 23, -38, 22, -115, -63, 42, 30, 8, -24, -1, 127, 68, -91, -77, 12, 0, 72, 13, -125, -11, 81, 70, -24, -112, 19, 19, 43, 17, 26, -54, -87, 60, 65, 85, -94, 0, 116, -35, -128, -91, 127, 127, -28, -92, -92, -12, 103, -60, -25, 127, -83, -97, 47, 87, -63, 27, 100, 6, -113, -54, 127, -58, 0, 56, -123, -54, 61, -32, 72, 58, -128, 72, 38, -116, -51, 108, 18, 7, 79, -128, 23, -1, -71, 31, 54, 86, -128, 13, 94, -61, -42, 21, 114, -53, -102, 1, 51, 106, -38, -35, 13, -128, 42, 25, -89, 127, -99, -21, 127, -18, -128, 15, -13, -32, 4, 51, 45, -128, 63, 110, -7, 9, -26, -39, -40, 63, -44, -128, 127, 71, -17, -40, -10, 14, -11, -63, -31, 123, -95, -34, 110, -58, -58, 69, 91, -64, -32, -48, 34, 19, -123, 75, -5, 49, -7, -36, 111, -88, 19, 52, 25, 29, -128, 63, 13, -24, 127, -24, -60, -100, -13, 17, 3, 72, 79, -62, -128, 52, 45, 46, 27, -41, -78, 65, -1, -79, 26, 74, 52, -128, -13, 85, 30, -1, -86, 88, 0, -124, 75, 97, -74, 20, 109, -42, -70, 43, -104, -11, 51, -46, 28, 85, -93, -43, 127, -92, -91, -10, -8, 120, -18, -25, 12, 18, 127, -82, -46, -36, 27, -20, 68, -13, -128, 127, 96, -66, -2, 37, -51, -128, -2, 127, -94, -86, 127, 19, 8, -6, 1, 31, -88, 26, -4, -72, 77, -40, -106, -1, 85, 66, -23, -38, 54, 8, -51, 5, -17, -47, 14, 93, -37, 10, 71, -91, -47, 11, -27, -31, -21, 127, 127, -115, 5, -9, -128, 51, 111, -106, 47, 0, 5, 12, -30, 54, 23, -49, -124, 15, 59, 41, 64, 54, -110, -8, -35, 38, -36, -91, 127, -69, -109, 127, 44, -110, -81, 102, 86, -14, 28, -28, -128, 40, 127, -7, -102, 19, -55, -28, -8, 14, 5, 62, 62, -97, 47, 34, -65, 11, -20, -97, 127, 48, -128, 6, 127, -46, -89, 72, -20, -53, 10, 14, -19, -29, 14, 75, -54, -29, 43, -94, 127, 39, -128, 48, 127, 40, -113, -74, 60, 20, 10, 8, -109, 62, 127, 15, -128, -78, 94, -4, 18, 65, 3, 26, -126, -127, 108, -22, -6, 108, -81, -34, 127, -51, -128, 127, -7, -103, 27, 24, 106, -5, 27, 24, -106, 37, 43, -55, -46, -41, -54, 127, -18, -39, 127, -128, -128, 73, 29, 45, -52, -6, 43, -125, 127, 3, -24, 127, -108, 29, -4, -128, 69, -9, 29, 127, -128, -68, 97, -57, 36, 41, -87, 56, 32, -121, 114, 43, -53, -9, -94, 90, 127, -94, 0, 70, -49, 4, 13, -115, 40, -21, -66, 65, -25, -1, -8, 6, 76, 43, -18, -45, -103, 127, -37, -63, 39, -106, -8, 127, 29, -110, 80, -28, 24, 71, -128, 23, 43, 29, 96, -128, 56, 18, -77, 28, -13, 96, 24, -95, -4, 11, 11, 76, -55, -128, 19, 127, -127, 7, 95, -95, 119, -61, -76, 127, -26, 1, -38, -128, 75, 21, -77, 92, 12, 28, 110, -128, -19, 127, -62, -29, -35, -1, 14, 66, 14, -128, 30, 79, 32, -107, 31, 127, -128, -8, 53, 44, -51, -11, 104, -23, 41, -128, -81, 95, -100, 0, 95, 63, -58, -109, 39, 64, 34, 47, -24, -100, -64, -25, 127, 113, -128, 19, 66, -77, 0, -58, -22, 103, 112, -115, -61, 127, -59, -128, 34, 39, -2, 127, -92, -17, 5, -46, 41, 46, -4, 22, -60, -63, -8, 87, 43, -128, 104, 74, 5, -128, 64, -26, -24, 127, -128, -51, 106, -3, -17, -56, -108, 24, 34, 0, -32, 12, 127, -2, -98, -12, 26, -1, 69, 11, -69, -75, 98, 24, -128, 114, 48, 30, 80, -128, 52, -18, -128, 127, 127, -11, -123, -113, 17, 70, 35, -59, 119, -27, -15, 8, -34, 3, 12, 27, 20, -60, -40, 117, -73, 4, -5, 20, 63, -112, -65, 83, 26, -62, 17, 22, -68, 53, 54, -52, -69, 96, 66, 38, -89, -95, 54, 34, 53, 60, -95, -71, 1, 59, 2, -60, 58, 2, -43, 89, 75, -120, 18, -81, 13, 127, -103, -18, 35, -3, -81, -27, 86, -7, 8, -35, 79, 51, -128, -11, 119, -96, 66, 76, -5, -93, -128, 58, 64, 9, -44, -39, 86, 115, -127, -54, 109, 0, -83, -35, 6, -6, 86, 48, 15, -68, -128, 103, 127, -106, -102, 72, 26, -44, -30, 30, 20, -10, 49, 82, -11, 31, -119, -72, 127, -53, -128, 41, 127, -71, 3, -41, -32, 79, 12, -19, -24, 103, -116, -28, 0, -21, 3, -1, 121, -72, 27, 127, -56, -85, 64, -24, -83, 105, 86, -128, -89, -41, 108, 13, -102, 110, -63, 91, -48, -1, 61, -66, 96, -48, -98, 62, 112, -105, -91, 45, 53, -74, -2, 2, 37, 19, -15, -13, -59, 80, 14, -3, 37, -69, 15, 121, -5, -10, 10, -14, 13, -115, -32, 78, -5, 51, -54, -35, -51, 51, -28, -25, 127, -79, 11, 1, -17, -13, -9, -45, -116, 14, 109, 66, -59, -31, 37, -25, -42, 55, -29, -56, 102, 81, 15, -62, -15, 6, -128, 127, 12, -128, 127, -48, 1, 108, -40, 14, -89, -40, 127, -59, -26, 40, 51, -97, 13, 82, -116, -29, 106, 36, -96, 48, -31, -39, -6, -75, 125, 46, -128, 127, 70, -38, -59, -74, 70, 95, -102, -7, 48, 27, -37, -128, 79, 127, -75, -98, 71, 0, 55, -56, 83, -51, -1, 44, -85, -13, -24, 37, -2, 29, -53, 116, -20, -106, 36, 56, -15, -59, 41, 38, -34, -26, 60, 38, -51, -9, 121, 9, -128, -11, 127, -128, -53, 127, -82, -102, -54, 93, 77, -58, -73, 69, 47, -88, -39, 52, 127, -105, 27, -3, -21, -15, -23, 36, -9, 109, 15, -42, -68, 81, -61, -97, 127, 64, -112, -76, -34, 28, -23, 14, 127, -108, -70, 18, 0, 31, 68, -40, -28, 86, -37, -52, 38, 122, -26, -128, 85, -8, 20, 10, -108, -34, 105, 32, -128, 2, 114, -32, -7, 85, 13, -54, 21, -65, -29, 13, -26, 36, -58, 127, 74, -63, -81, -34, 64, 45, 19, -45, -105, 45, 123, -66, 8, 35, -27, 39, 31, -109, 51, 12, -17, 59, -35, -3, 1, -71, 17, -32, -31, -8, -83, 52, 86, -19, 14, -44, 70, 28, -124, 127, 65, -128, -63, 76, 66, -96, -62, 106, -9, -56, 125, 3, -128, 127, -35, 18, 22, -7, -15, -41, 127, -128, 45, 57, -124, 51, 19, -56, 44, 116, -108, -31, -40, 24, 3, 0, 110, -65, -86, 103, 96, -128, -73, 109, 122, -114, -30, 0, -115, 110, 107, 11, -6, -9, -79, -87, 8, 96, 40, -128, 34, 127, -28, -8, -41, 14, 18, -115, -43, 127, -53, 24, 127, -128, -19, 89, -17, -94, 56, 88, -128, 22, 100, 0, 5, -128, -75, 127, 85, -40, -124, -26, 90, 39, -41, -128, 64, 127, -100, 19, 66, -114, 76, -3, -17, 46, -94, -28, 127, -43, -124, 7, -57, 127, -31, -78, 127, -117, -59, 105, 34, -4, -117, -15, 40, -5, 36, -86, -51, 127, 74, 9, -128, 4, 8, 37, 6, -78, 45, -71, 78, 66, -107, 56, 43, -97, 8, 25, -19, 127, -64, -127, 127, -28, 44, -62, 12, 69, -128, -1, -21, 127, 127, -128, -59, 127, 52, -63, -66, -90, 100, -37, -12, -11, 25, 23, -105, 32, 13, 102, -72, -40, 127, 9, -34, 1, -7, -27, 39, 32, -78, 49, -1, -77, -75, -54, 61, 127, 27, -11, -106, -55, 127, 21, -69, -20, 52, 4, 1, -87, -76, 121, 51, -114, -13, 57, -110, -15, 35, -59, -14, 127, -54, -5, 78, -128, 123, 127, -128, 5, 120, -95, -55, 86, -66, 66, 59, -128, 120, 24, -89, 37, -34, -26, 81, 102, -13, 6, -110, 27, 127, -128, -9, 115, -128, 38, 127, -26, -27, -3, 6, -92, -88, 109, 127, -128, 22, 10, -125, 98, 8, -26, 91, -30, -26, 10, -79, 3, -17, 9, -7, 81, 61, -24, 1, -41, 40, -47, -23, 14, -41, -44, 81, 54, -128, 41, 89, 39, 8, -4, -24, -128, 13, 30, 36, -52, 13, 127, -97, 31, -45, -61, 104, 18, -54, -78, -12, 127, 18, -39, -30, -15, 95, 44, -128, 10, 75, -66, 82, -104, -22, 25, -74, 127, 17, -44, 115, -128, -49, 61, -128, 66, 127, -31, -68, -90, 80, 98, -128, -41, 66, -18, 126, -34, -121, 11, -54, 117, 95, -15, 44, -89, -128, 14, 19, 35, 127, -98, -46, 102, -72, 44, -31, -66, 18, 54, 25, -92, -25, 79, 11, -3, 97, -62, 6, -29, -82, 127, 76, -128, -24, 127, -76, -14, 97, -25, -128, 68, 106, -128, -9, 43, 6, 105, -28, -128, 13, 2, -68, 127, 38, -25, -27, -13, -43, -51, 114, 56, -108, 11, 104, 45, -56, -119, 75, 9, 13, 121, -114, -58, 121, 17, -21, -30, -22, -48, 31, -47, -74, 127, 79, -128, -24, 59, -49, 76, 1, -89, -51, 89, 63, 49, -60, 47, -40, -128, 63, 127, -93, -43, 127, -128, 22, 85, 5, -5, -128, 46, 100, -34, 1, -3, 6, -68, 27, 127, 1, -128, 56, 127, -82, -37, 29, -99, -20, 127, -123, 40, 125, -128, 28, 41, -97, 3, 127, -93, -34, 127, -57, -91, -4, -49, 63, 127, -125, -61, 104, 68, -43, -35, 51, -87, -65, 48, 9, -89, -20, 121, -54, -113, 127, 115, -77, -109, -26, 64, -49, 127, 7, -59, 29, -32, 112, -103, -64, 127, 14, -128, 102, 11, -128, 126, 82, -69, -15, -87, 37, 109, -6, -23, 23, -23, -54, -47, 24, 70, -26, 9, -2, 24, -59, 32, -9, 20, 115, -86, 44, -57, -8, 102, -76, 25, 26, -128, -36, 127, -78, -1, 80, -44, 3, -78, -58, 108, 19, -36, -18, 37, -36, -14, 55, -91, 12, 47, -39, -59, 10, -30, 83, -41, 80, 0, -8, 100, -128, -8, 44, 21, -20, -53, -12, 127, 12, -77, 91, -117, -70, 40, 77, 76, -128, -46, 127, -10, 0, -55, -26, 0, -79, 49, -36, -4, 57, -46, 64, 106, -66, -44, -55, 109, 42, -71, 54, 95, -122, -38, -10, -34, 127, 63, -128, 23, 44, -128, 60, 7, -15, -5, -19, 92, 0, -57, 80, 46, -75, -12, -30, 53, 83, -93, 8, -61, 64, 57, -128, 127, 127, -128, -45, 126, 55, -19, -42, -83, 53, -29, -65, 35, -68, 103, 82, -73, 74, 0, -128, 4, 127, -19, -128, 45, 82, 17, -17, -44, 77, 17, -98, 59, 7, 35, -9, -82, 59, -89, 31, 68, -108, -34, 71, 7, 61, -42, -20, 127, -77, 27, -63, -115, 127, -55, -72, 91, 6, -100, 53, 77, -80, -12, -51, -24, -7, 100, 41, 6, 43, -83, -108, 127, 22, -42, -13, -99, 111, 106, 22, -121, -48, 127, -52, -78, 127, -96, -128, 127, -42, 69, 0, -75, 51, -81, 88, -6, 51, -32, -128, 102, 37, -64, 3, 70, 76, -59, 1, 24, -98, 30, 57, 35, -11, -128, 1, 95, -78, 18, 19, -73, 81, -10, 39, 83, -56, -72, 122, -15, -99, -24, 53, 121, -100, -96, 6, 127, -13, 6, 0, -69, 27, 64, -35, -15, 108, -44, -79, -115, -19, 98, -39, 22, 81, 27, -56, -126, 0, 34, 20, 49, -35, 110, -29, -91, 2, -17, 74, -5, -15, 80, -81, 17, 127, -114, 30, 58, -109, -78, 105, 20, -24, 97, -120, -89, 127, -15, -64, 91, 11, -12, -59, 20, 87, -82, -73, 57, 82, -8, -107, -79, 77, -34, 126, -18, -100, 127, 4, 11, -128, -31, 35, 43, 20, -73, -47, 121, 93, -123, 53, -40, -128, 127, 126, -48, -90, -95, 53, -39, 57, 91, -120, -61, 100, -5, -72, -1, 114, 120, -38, 17, -75, -128, 66, 105, -76, 15, 28, 56, -79, -100, 22, -11, 9, 121, 122, -90, -128, -9, 65, 74, 37, -21, -128, -44, 127, -76, -53, 125, -107, -46, 111, -23, -8, -52, 91, 93, -46, -32, -32, 70, 6, -17, -100, -128, 127, -9, -60, 127, -26, -128, 94, 17, -15, 95, -32, -4, -128, -42, 88, -75, 60, 127, -66, -110, -43, 29, 127, 55, -8, -49, -23, 41, -98, 32, 92, -128, -123, 76, -11, 13, 74, 38, 63, -104, -15, 74, -128, 52, -8, -85, 127, 41, -85, -90, 127, 12, -64, 110, -81, -34, 63, -99, 12, -29, -55, 79, -12, -27, 114, -30, 13, 25, -128, 83, 76, 31, -75, -20, 74, -81, -73, 52, -29, -3, 127, -98, -128, 126, -22, -18, 51, 8, 108, -128, 27, 41, -89, 7, 21, 19, -15, 32, 9, 65, -83, -54, 99, 31, -80, -4, -43, 41, 3, -66, 73, -71, 34, 81, 9, 42, -98, -89, 95, -26, -62, 83, -10, 36, 43, 41, -107, -119, 76, 99, -97, 3, 38, 8, 28, -35, -1, -8, 3, -28, 112, 27, -69, -14, -39, -14, -3, 23, 44, 52, -8, 8, -25, -128, 85, 23, -128, 127, 49, -80, 45, -2, -88, 91, 0, -52, 48, 4, -66, 54, 6, -128, 93, 95, -7, 51, -115, 31, 64, -68, 115, -128, -9, 53, -99, 35, 44, -29, -56, 106, 69, -17, -93, 24, 62, -87, -29, 80, 100, -104, -56, 114, -62, 29, 13, -26, 71, -99, 36, -51, -119, 121, -20, 20, 127, -89, -102, -7, 72, 20, -98, 0, 9, -32, 127, 28, -88, -18, -36, 18, 31, 94, -102, 18, 114, -86, 25, -39, 53, 13, -86, -29, -85, 93, 127, 1, 35, -127, -128, 114, 52, -100, 73, 56, -103, 51, 91, -11, 22, -103, -128, 59, 127, -56, -113, 80, 53, 54, 34, -51, -76, -44, 76, -15, 41, 55, -128, 83, 82, -128, 4, -47, 3, 34, -19, 83, 74, -85, -73, 104, -34, -28, -27, -68, 110, 0, 6, 5, -92, 45, 111, -22, 0, -6, 1, 68, -128, -111, 121, 102, -53, -108, 102, -61, -65, 76, 28, 2, -6, -12, -77, -30, 117, 39, -102, 30, 83, -107, 41, -13, -53, 127, -35, -22, -46, 13, 13, -27, 86, -60, -68, 35, 27, -10, -19, -6, -117, 20, 127, 20, 1, -82, -128, 124, 110, -75, -36, 10, 52, -43, 2, 29, -82, 15, -27, 70, -13, -6, 73, -115, -19, -26, 81, 127, -43, -91, -36, 29, 108, -78, -91, 114, -7, -63, 46, -80, 95, -37, -59, 127, -79, -21, -49, 38, 127, -83, -49, -24, -83, 127, 5, -109, -3, -57, 51, 110, -3, 8, -12, -79, 122, 74, -128, -27, 17, 40, 78, -122, 49, 7, 25, -35, -7, -29, 8, 122, -108, -43, 61, 34, -96, 77, 108, -128, 56, -41, 4, 42, -26, -13, -35, 127, -128, 42, 54, -128, 80, 96, -37, -68, -36, -5, 55, 102, -42, -89, 40, 41, 45, -94, -70, -9, -10, 5, 40, 2, -24, 39, 49, -58, 30, 13, 36, 87, -128, -89, 127, 82, 0, -49, -128, -28, 100, 74, 28, 90, -128, -77, 127, 26, -21, 27, 9, -4, -124, -128, 127, -7, -95, 52, -60, 115, 55, -128, 19, 108, -89, -27, 11, 108, 68, -128, 114, -30, -47, 127, -128, 11, 48, -21, 71, -128, 54, 48, -2, 76, -89, 36, -120, 48, 40, -128, 127, 59, -127, -15, -10, -19, 97, -4, -64, -22, 66, 1, -47, 54, -48, 23, 17, 9, 0, 53, 71, -128, -38, 75, 85, 59, -123, 12, 97, -79, -125, 75, -12, -55, 19, -49, 112, 73, -57, 36, 78, -128, -108, 36, 58, -7, 20, 74, -6, 46, -29, -119, 97, 72, -49, 24, -18, -128, 44, 52, -53, 106, -106, -17, 44, -119, 119, 108, -12, -102, 0, 71, -97, 42, 66, -45, 62, -74, -121, 98, -59, 11, 125, 31, -73, -71, 62, 62, -19, -89, -30, -28, -13, 25, 103, -12, -61, 59, -49, -73, 127, -94, 7, 49, -45, 69, 11, 9, -4, -73, -112, 127, 119, -128, 23, 46, -61, 79, -73, -31, -40, 58, 83, -61, -70, 3, 117, 46, -128, -78, 18, -14, 27, -17, 45, -24, 58, 49, -9, 47, -19, -90, -3, 105, -80, 13, -31, -94, 62, 57, 18, 14, -38, -80, 127, 31, -83, 114, -108, 17, -8, -116, 127, -28, -97, 35, -10, -49, 93, -25, 4, 65, -110, 0, 127, -3, -29, 100, -71, -125, -25, 127, 35, -108, 98, -13, -36, 45, -125, 94, 14, -127, 12, -15, 43, 61, -20, 26, 43, -128, 44, 41, -93, 119, 30, -113, -34, 44, -44, 56, 65, -75, 45, -87, 49, 95, -94, 49, -83, 18, 96, -57, -111, 77, 110, -78, -18, -60, -6, -10, 11, -1, 0, 127, -82, -111, 30, 40, 79, -18, -57, -38, 102, 127, -128, -2, 38, 6, 0, -38, 57, -88, -90, 127, -17, -128, 70, 119, -36, -128, -72, 127, 11, -74, 119, -65, -1, 102, 5, -83, -62, -48, 69, 32, -102, -14, -5, 127, -51, 3, 92, 11, -90, 7, 127, -105, -120, 30, 23, 2, 47, -49, -17, 61, 92, -99, -128, 127, -34, 57, 4, -86, 6, 41, 127, -128, 58, -32, -128, 12, 127, 83, 20, -120, -54, 127, -70, 13, -32, 0, 6, 21, -55, -7, 114, -128, -97, 123, 127, -128, -10, 127, -38, -14, 28, -54, -115, 56, 75, -122, 68, 7, 5, 77, -110, -11, 22, 57, -45, 0, 53, -31, 13, 0, -5, -92, 49, 76, -128, 3, 127, 6, -46, -47, 35, -49, 55, 104, -128, -48, 127, 24, -47, 25, -47, -112, -21, 127, -99, -56, 127, -44, -58, -5, 3, -99, 103, 12, -49, 125, 5, -72, -17, -1, -114, -8, 107, 127, -128, -35, 107, -128, 37, 22, 78, -54, -82, 92, -105, 56, -12, 73, 4, -64, 66, -26, 61, -69, 29, 38, -127, 46, 125, 5, 0, 41, -128, -38, 127, -111, -75, 60, -58, 103, 81, -128, 93, -11, -76, -13, 11, 99, 10, 48, -128, -68, 27, 87, 46, -128, -53, 111, 92, -125, -28, 127, -120, 5, 58, 24, 78, -26, -73, -128, 121, -26, -104, 127, -65, 7, 110, -22, -55, -23, 32, -25, 53, 55, -96, -44, -77, 45, 26, -11, 104, -8, -71, 27, -12, -9, 83, -122, 10, -24, -52, 91, -83, 70, 25, -102, 66, 127, -92, -128, 126, 95, -13, -17, 3, -65, -93, 88, 125, -73, -81, 83, -80, 43, 66, -88, 70, -74, 27, 31, -89, -24, 91, 14, 0, 111, -58, -90, 66, 41, -82, -2, -9, -53, -49, 127, 26, -128, 91, -31, -28, 127, 6, -73, 2, 76, 56, -128, -128, 90, 61, -81, 63, -42, -22, 57, 37, 103, -42, -53, -5, -81, -88, 127, 11, -128, 111, 39, -70, -30, 18, 85, 76, 56, -128, -71, 127, -128, 0, -6, -28, 55, -82, 31, -18, 78, 79, -128, 35, 38, 2, -9, -74, 127, -97, -52, 127, 3, -128, -75, 127, -5, 3, 86, -99, -107, 20, 45, -38, -18, 11, 121, -10, -35, -46, 13, 37, -4, 96, -127, -107, 106, 15, 6, 12, -36, -18, 7, -22, -24, 83, 103, 0, -75, 43, -97, 12, 24, -78, 127, -42, -29, 82, -13, -38, -128, 10, 127, 34, -124, 36, 107, -27, -105, -31, -9, 17, 99, -45, 26, -88, -108, 127, 65, 4, -55, 15, 6, -28, -29, -17, -27, -59, 76, -69, 65, 73, -64, 64, -79, 41, 91, -128, 24, 127, 0, -128, 14, 102, -30, 2, -18, 82, -61, -94, 88, 74, -83, -83, 56, 44, 44, 21, -128, -62, 127, 38, 3, -73, -46, -36, -24, 11, 8, -7, -26, 20, -30, 127, 77, -30, -20, -86, 57, 71, 3, -49, 3, -77, 62, 14, -25, 127, -128, 43, 30, -31, 113, -128, -56, 35, -25, 68, 6, -19, 54, -26, -8, 49, -49, -76, 24, 81, 20, -113, 10, 26, 31, -28, -39, 87, -10, -29, 4, 39, -34, 41, 38, -105, -100, 127, 76, -128, 15, 85, 70, -128, -82, 66, 77, 11, -15, -56, -51, 10, -10, 106, 30, -128, -68, -2, 109, 64, -38, -39, -83, 127, -46, -34, 49, -128, 103, 90, -46, -81, 34, 29, -55, 96, 90, -128, -36, 79, -31, 62, 45, -11, 9, -107, 46, 81, -115, 2, -35, 42, 103, -122, 6, 100, -128, 25, 127, -69, -38, -87, 44, 127, -103, 22, 75, -128, -68, 7, 79, 44, 63, -31, -113, 74, 53, -73, -21, -52, 88, 88, -14, 32, -128, 36, 97, -128, 59, 19, 19, -26, -56, 62, 78, 62, -112, -24, 97, -39, -23, 18, -128, 45, 127, -71, -71, 13, 52, 48, -43, -17, -12, -14, -21, 4, -19, 47, 38, 29, -85, -125, 127, 0, -69, 120, -88, -128, 102, -21, 20, 37, -35, 100, -116, -36, 36, -28, 123, 82, -128, -65, 66, 44, -126, 56, 41, -128, 99, 87, -114, 15, -6, -98, 21, 121, -18, -93, 127, 34, -82, 25, -77, -74, 95, -31, 39, 88, -29, 0, 21, -128, -59, 61, 73, -1, -74, -68, 94, -19, -8, 127, -53, 20, -128, 12, 127, -128, -43, 76, 81, 52, -93, -128, -14, 127, 13, -128, 104, -13, 23, 80, -128, -41, 127, -65, -37, 69, -128, 54, 12, 85, 21, -128, 112, 43, 19, 7, -60, 3, -102, 69, 24, -32, 76, 2, -29, -96, 63, 24, -100, 85, 74, -48, 37, 26, -71, -6, 59, 22, -128, -68, 114, 22, -61, -7, 115, -52, 5, 52, -82, 127, -117, -9, 85, -32, -8, 19, 90, -128, -97, -3, 98, 123, -59, -22, 0, -90, -22, 31, 95, -28, -38, 17, 0, 78, -1, -41, -119, 10, 127, -18, -56, -98, 15, -2, 26, 127, -128, -24, 51, -119, 119, 127, -128, -87, 127, 3, -26, 61, 66, -94, -113, 34, 77, 71, -83, -64, 29, -9, -56, -22, 127, 27, -124, -7, 65, -65, -39, 87, 55, -31, 0, 14, -71, 36, 108, -128, -102, 82, 117, -79, 0, -2, -43, 109, -119, -78, 10, 73, 61, -89, 87, 32, -17, -46, 31, 42, -111, 24, -53, -44, 127, 91, -35, -79, -17, 74, -27, -126, -21, 96, -9, -66, 105, -55, 9, 127, -128, -128, 58, 110, -41, -51, 2, -55, 97, -5, -40, 127, -29, -62, -31, -28, 73, -104, 91, 10, -18, 57, -109, -42, 123, 63, -116, 30, 49, -74, -21, 107, -64, 35, 20, -62, -21, -7, 69, 26, 17, -128, 56, -5, -38, 127, -37, -128, 110, 42, -128, 89, 69, -69, 35, 32, -128, -36, 32, 57, 34, 9, -30, 13, 35, -4, -54, 19, -19, 21, 39, 0, -76, -125, 127, 64, -128, -31, 127, -86, 17, 24, -128, 97, 110, 42, -103, 3, -4, -62, 55, 36, -59, 28, 43, -17, 17, -4, -3, 1, 47, -128, 11, 125, -90, 9, 6, -7, -27, -76, 127, -55, -77, 127, 31, -126, 40, -30, -116, 8, 69, 88, 0, 40, -44, -106, 63, -24, -104, 70, -51, 107, 66, -40, 35, 17, -3, -128, 19, 123, -31, -31, -78, -65, 82, 112, -8, -69, -97, 71, 80, -35, 0, -64, 11, 110, 12, -115, -94, 105, 95, -128, 58, -24, 37, 83, -128, 43, 97, 15, -30, -75, -8, 48, 3, 68, 2, -128, 5, 62, 65, 79, -128, -78, 17, 77, -12, 40, -43, -102, 127, 14, -27, -36, 34, 40, -128, 86, 35, -69, 96, 6, -113, -96, 61, 85, -68, 37, 117, -73, -57, 38, 8, 7, -86, 37, 78, -92, 76, -1, 26, 20, -128, 38, -12, -87, 46, 9, -41, 55, 124, 47, -128, 15, 127, -80, -56, -86, 1, 28, 3, 93, 22, 48, -99, -18, 76, -18, -79, -35, 24, -45, -41, 54, 127, -99, 3, -5, -82, 127, 37, -113, 2, 127, -108, -43, 66, -5, 19, 23, 55, -128, -31, 119, -89, -125, 111, -40, 19, 127, -81, -110, -52, 69, 127, -128, 17, 121, -128, -28, 41, 86, 36, -128, 43, 121, -12, -85, -30, 45, -54, -3, 64, 103, -119, 23, -28, -40, 127, -19, -21, -63, -90, -66, -22, 127, -26, -128, 127, 21, -79, 127, 102, -15, -128, 0, 107, 6, -91, -104, 63, 8, 75, -63, -68, 127, 102, -104, -45, 120, -83, -60, 29, -10, 18, 5, -6, -6, 29, -103, 21, 127, -128, -18, 127, -128, -20, 41, 63, 30, -63, -69, 83, 2, -128, 47, -27, -17, 97, 110, -93, -126, 55, 91, 44, -122, -44, 40, 66, -59, -52, 87, 73, 4, -128, 45, 54, 30, -108, -23, 68, -15, 95, -81, 34, -44, -27, 0, -60, 105, -112, 46, 120, -62, -15, -18, 10, 79, 14, -79, -125, -29, 127, 93, -30, -121, -10, 66, -125, 81, 0, -51, 96, -93, -85, 99, 22, 36, 55, 0, -59, -17, 73, -127, -30, 20, 49, -25, -78, 76, 52, -57, 40, 58, -110, 14, 92, 66, -128, 14, 127, -128, 0, 14, -44, 59, 70, 10, -66, -21, 11, 65, -40, -128, 127, 70, -114, -1, 48, -12, 69, -94, -26, 103, -71, 83, -81, -121, 127, -41, -107, 74, 6, 38, 44, -4, -64, -30, 11, 27, 93, 17, -59, -128, 119, 30, -54, -1, 35, -10, -7, 98, -105, 0, -24, 61, 36, -99, -22, -32, 58, 14, -2, 98, -109, -104, 99, -14, 14, 66, 43, -53, -61, -13, 7, 12, 27, -53, 17, 58, -62, 44, -70, 71, -1, -83, 127, 2, 4, 59, 1, -99, -75, 43, -31, -21, 90, 22, -5, -57, -55, 44, 46, 32, -8, 47, 77, -128, 39, 85, -116, -24, 94, 39, -128, 103, 127, -68, -53, -9, 35, -82, 53, 109, -83, 53, -75, -128, 82, 76, -49, 24, -75, 40, 46, -81, 125, -100, -24, 116, -9, -110, -91, 95, 82, -96, 6, 39, 31, 94, 22, -91, -128, 122, -17, -20, 127, -124, 65, -21, 1, 8, -31, 127, -128, -126, 71, 127, -43, -128, 65, 127, -114, -27, 45, -24, 59, 3, 45, -71, -46, 76, -8, 2, -37, 18, 9, -90, -56, 43, 51, 89, 44, -128, 54, 86, -81, -66, 34, 65, -31, -92, 28, 49, 21, 69, -128, -70, 117, -122, 59, 25, -35, 44, 29, -40, -120, 49, 26, -26, 48, 109, -98, -55, 13, -38, 3, 90, 78, -128, 14, 48, -58, 38, -85, 10, 76, -59, 127, -41, -128, 127, -13, -128, 39, 25, -20, 69, 32, 37, -121, -63, 127, -64, 69, -66, -56, 61, 29, 15, -90, 43, 32, 38, 34, -20, -109, -77, 127, -28, -112, 58, -73, 73, 66, -73, 93, 74, -128, -19, 113, -94, -85, 44, 78, -64, -10, 15, 3, 17, 1, 96, 51, -124, -10, 91, 9, 63, -128, 23, 36, -99, 37, -24, -27, 69, 122, -128, -36, 127, 31, -128, 63, 127, -113, -49, 69, 54, -44, -86, -77, 0, -21, 127, 22, -38, 69, -112, 26, 83, -128, 36, 127, -128, 8, 127, -32, -68, 40, -41, -104, 79, -2, -42, -10, 79, 86, -128, -6, 48, -65, 65, 4, -51, 1, 68, -62, -112, -34, 123, 116, -128, 5, 99, -73, 4, 48, -62, -57, 62, 53, 21, -54, -91, -18, 127, -12, -128, 127, 121, -107, -35, 37, -62, -85, 48, -21, 14, 82, -62, -15, 15, -35, 127, 72, -77, -17, -62, 55, 65, -6, -44, -94, 127, 4, -115, 71, -5, -47, 63, -68, 79, -20, -20, 13, -128, 127, -56, -85, 104, -112, 82, 71, -116, 60, -44, 39, -4, -96, 89, 68, -106, 11, 127, 18, -128, -104, 95, 6, 36, -75, -12, 105, -89, -35, 83, 0, -52, 38, 98, 2, -42, 22, -113, 75, 35, -128, 112, -5, -19, -32, 72, 54, -30, 70, -77, -128, -64, 127, 23, -30, -90, 55, 62, -128, 17, 115, 10, -44, -4, -36, -35, 111, 127, -128, 31, -19, -69, 95, -14, -94, 69, 49, -38, 70, -62, -105, 96, 55, -119, -21, 26, -12, -6, 62, -1, 4, -17, 53, -51, -14, 10, -80, 93, 108, -12, -75, -57, -38, -10, 90, 12, 57, -56, 19, 116, -117, -48, -8, 127, -25, -32, -26, -32, 127, -11, 0, -52, 13, 43, -96, -2, 19, 44, -110, -12, 37, -27, 79, -44, -2, -30, 11, 43, -81, 29, 127, -14, -29, -38, -26, -11, -104, 109, 100, 32, -61, -47, 21, -40, -35, 121, -49, -128, 127, -2, -58, 127, 1, -128, -21, 5, -13, 127, 4, -64, 6, -14, -35, -54, 108, 87, -111, 36, 32, -128, 76, 126, -19, -98, -60, -10, -8, 52, -56, 126, 42, -88, 127, -128, 3, 68, -128, 25, -12, 73, 102, -12, -99, -83, -22, -23, 127, 49, -128, 14, 86, 77, -54, -75, -14, 43, 62, -64, 89, 32, -99, -18, -10, 1, 39, -45, 41, 91, -30, -128, 18, 76, 15, 68, -51, 24, -117, -35, 80, -128, 127, 123, -28, -87, -97, -38, 113, 110, -109, 48, -43, 24, -17, -43, 24, -13, 127, -128, -65, 104, -66, -88, 127, 127, -29, -52, -29, 81, -94, -128, 127, -12, -35, 127, -94, -128, 113, 13, -27, 36, -125, -22, 28, 19, 83, 8, 40, 14, -83, 5, -103, 48, 59, 43, 22, -120, 32, -1, -64, 97, 15, -116, 127, 7, -128, 40, 63, -83, 64, 34, -79, 126, -37, -18, -15, -104, 35, -7, 73, 100, -45, 2, -12, -128, 52, 127, -66, -107, -20, 102, -54, -31, 127, 26, 7, -128, -78, 73, -31, -54, 75, 110, -128, -104, 97, 13, -57, 92, 0, 46, -6, -1, 43, -56, 88, -105, -32, 26, -52, 95, 85, -74, -98, 109, -8, -85, -61, 75, 127, -100, -128, 63, 14, -106, 110, 72, -97, 83, -35, -54, 121, -40, -23, -23, -47, 32, 34, 68, 15, 12, 1, -47, -21, -90, 32, 127, -29, -36, 48, -40, -128, 109, -21, -108, 0, 56, 127, -104, -52, 114, 59, -128, -66, 42, 1, 34, 30, 68, -59, -100, 121, -56, -128, 72, 11, 81, -29, 25, 73, -128, -8, 127, -98, -19, 20, -91, 34, 127, -10, -27, 97, -128, 74, -18, -86, 70, 18, -22, -45, -35, 72, 35, -119, 121, 59, -71, 1, 71, -17, -112, -47, -19, -3, 14, 110, -22, -78, 127, 104, -62, -46, 12, 31, -21, 1, -21, -128, 29, 114, -35, -6, -5, 2, 91, -85, -82, 59, -80, -2, 13, -29, 98, -45, -36, 107, 58, -70, 55, 34, -115, 31, -10, -91, 37, 127, 55, 8, -128, -59, 125, -6, -74, -63, 44, -13, 13, 110, 0, -30, -88, 21, 122, -38, 7, -76, -77, 68, 49, -61, 75, 117, -39, -93, -124, 38, 38, -58, 20, 37, 30, 106, 24, -13, -116, -114, 127, 38, -9, 9, -128, -54, 0, 127, 58, -31, 58, 8, -123, -79, 127, -56, -128, 127, 3, -77, -43, 52, 47, -66, 82, 107, -124, -37, 98, -87, 36, 31, -3, 53, -128, -128, 127, 2, 0, 56, -128, 103, 29, -105, 21, -9, 34, 63, -91, 47, 127, -128, -54, 25, 17, 23, -82, 94, 127, 8, -128, 12, 80, -128, 38, 96, -96, -38, 127, -102, -12, 127, -8, -128, -97, 18, 6, 86, 38, -52, -24, 21, -1, 66, 2, 52, -110, -40, 127, -128, -20, 127, 30, -128, -113, 74, 115, -25, -128, 83, 63, 11, 40, -87, -123, 102, 76, -117, -4, 122, 8, -39, -14, -128, 34, 127, 59, -81, -47, 44, -18, -78, 41, 21, -57, 75, 91, -100, -100, -19, -47, 125, 127, -8, -128, 59, 81, -79, -26, -106, 53, 127, 4, -5, 32, -124, -4, 94, -12, -59, -39, -24, 57, -41, 3, 30, -128, 105, 89, -102, 41, 73, -128, 34, 65, -106, 91, -69, 14, 127, -128, -85, 127, 54, -102, 7, -23, -105, 113, -69, 35, 28, -85, 86, -5, -82, 86, 26, 14, -20, -30, 51, 15, 51, -115, -62, -9, -60, 63, 3, -71, 83, 59, 85, -58, 2, 81, -80, -66, -29, 88, -79, 9, 1, -25, 127, -91, -97, 69, -73, 77, -5, -11, 88, 51, -128, 30, 34, -128, 92, 6, -71, 127, 59, 39, -88, -82, 127, -14, 32, -94, -106, 127, 57, -110, -29, 61, -4, 17, 86, -43, -105, 125, -66, -10, 127, -128, 17, 127, -128, -86, -7, 2, -2, 61, 35, -85, -23, 127, 88, -32, 31, 8, -45, -56, -95, 82, 127, -107, -53, 53, 41, 20, -18, -128, 54, 115, -128, 70, 61, -89, -60, 25, 96, -69, -104, 127, 25, -128, 112, -36, -127, 112, 127, 10, -128, -109, 127, -25, -14, 39, 34, 58, -123, 21, 80, -71, -83, 127, -49, -10, 56, -108, 51, -69, 22, 92, 29, 41, -12, -54, 6, 78, -128, -2, 95, -128, 75, -1, -105, 48, 39, -35, -113, 116, 127, -38, -112, -102, 115, 28, -115, -45, 121, 77, -120, -13, 20, -44, -4, 127, 83, -128, 59, 127, -128, -27, 89, -122, -57, 127, 73, -19, -87, 0, 124, -128, -27, 127, -61, -105, 15, 19, -4, 96, 89, -93, -113, 115, 41, -128, 126, -62, -88, 127, -112, -52, 108, -51, 9, 39, -63, -61, 26, 6, 87, 107, -104, -98, 89, 29, -57, 63, 42, -34, -1, -13, -125, 80, 57, -76, -11, -38, 56, 82, -92, -6, 20, 21, -63, 35, 59, -128, 127, 36, -120, 91, -43, 5, -18, -128, 46, 78, 112, -107, -96, 117, 32, -38, 6, -90, 80, 127, -128, -17, 30, 6, -71, 61, 21, -128, 95, 45, -66, 60, -100, 46, 103, -128, 51, 49, -47, -104, -12, 71, -53, 39, 127, 10, -128, -36, 127, -87, -79, 26, 54, 102, -9, 13, 1, -128, -70, 64, 65, 51, -108, 12, 88, -2, -90, -44, 57, 20, 1, 3, 85, -22, -119, 85, -9, -85, 46, -75, 28, 108, -55, -73, 59, -25, -52, 32, -1, 27, 53, 100, -121, -9, 103, -27, -19, 14, -40, -128, 45, 116, 39, -64, -52, -35, -11, 99, 30, -8, 55, -103, -46, 6, -17, 127, -62, -34, -4, -19, -17, 55, 73, -128, 77, -9, -116, 24, 127, -9, -128, 54, -39, -81, 127, 53, -122, -18, -29, 104, 119, -18, 37, -128, 27, 46, -128, 12, -19, 3, 127, -42, -95, 29, 15, 127, -25, -68, -4, -42, 117, 11, -27, 72, -41, -38, -58, 30, 85, -94, -22, 52, -69, -19, 124, -81, 0, 127, -116, 11, 0, -123, -24, 61, 52, -10, -5, 70, -90, -4, 21, 29, 38, -128, 111, 127, -44, -128, 41, 41, -44, 15, -123, 86, 127, -4, -128, -7, 127, -78, 2, -62, -1, 119, -6, -107, -41, 30, -72, 69, -18, -39, 96, -14, -7, 7, -5, -51, 61, -7, 1, 12, -26, 100, -102, -29, 98, -62, -40, 31, 96, -86, -20, 89, 39, -32, -11, -7, 0, -48, -128, 127, 52, -66, -27, 88, -70, -27, 36, -39, 127, -10, 5, -39, -59, -55, -62, 10, 43, 42, 40, -55, 1, 9, 39, 34, -20, 58, -128, -9, 127, -128, -19, 37, -9, 127, -108, -30, 96, -70, -39, 59, -36, -27, -6, 65, 65, -109, 75, 98, -39, -45, -102, -36, 127, -106, 8, 127, -45, -117, -61, 127, -93, 69, 121, -68, 3, 52, -72, -82, -10, 83, -68, -36, 49, -68, 26, 80, 43, -98, 39, 10, 12, 81, -26, -23, 15, 8, -74, -19, 45, 52, -125, 1, 110, -1, -35, -69, 57, 85, -128, -128, 127, -68, -21, 127, -105, -128, 82, 127, -72, -73, -3, -14, -22, 127, 107, -12, -17, -116, 6, 34, -96, 82, -8, 23, 74, -41, -13, -52, 53, -18, 1, 0, -42, 12, -35, 47, 38, -128, 0, 127, -76, -5, -46, -54, 113, 62, -35, -92, -5, -60, 104, 42, 15, -62, -78, 92, 87, -99, -128, 127, 74, -128, -31, 40, 22, 116, -104, -116, 127, 75, -128, -52, 75, -42, 76, -7, -121, 46, 58, 18, -15, -31, 107, -9, -89, 20, 89, -6, -76, -18, -43, 7, -3, 74, 4, 55, -9, -57, -34, -28, 27, -24, 69, 59, -31, -49, 58, 25, -9, -74, 52, 127, -117, 4, -43, 22, 13, -128, 25, 97, -2, -58, 103, -17, 43, -55, -108, 40, 44, 7, -27, 70, -26, 72, -71, -14, 10, -5, 8, -30, 104, 49, -36, -128, 60, 77, 11, 30, -24, -120, -55, 127, 1, -128, 4, 52, -45, 45, 52, -3, 43, 52, -96, -128, 127, -7, 5, 96, 17, -128, -80, 127, 60, 27, -39, -36, -42, 11, 0, -95, 51, 127, -124, -127, 127, 21, -77, -62, 74, 127, -77, -34, 21, 18, 14, -44, -128, 61, 58, -128, 76, 123, -24, -20, 2, -24, -55, -34, -1, -86, 70, 8, 14, 127, -128, 36, -31, -11, 127, -128, -3, 115, -128, 24, 127, -128, -46, 127, 46, 4, -128, -25, 127, -128, -36, 127, 12, -97, -76, 22, -25, 127, 25, -128, 80, 127, -128, -128, 127, -22, -87, 120, 61, -52, -52, 22, -19, 78, -5, -113, 85, 49, -128, 36, 88, 0, -17, -79, 98, 48, -62, -86, 42, -35, -55, 85, 64, -10, -56, 36, -30, 74, -45, -111, 27, 60, 57, 2, -19, -99, -66, 35, 108, -24, -121, 17, 127, 3, -68, 111, -98, -87, -5, 108, 22, -66, 32, -62, -32, -54, 127, 119, -128, -55, 13, 9, 127, 64, -128, -52, 127, -66, -19, 78, -86, 39, 85, -72, -107, 60, 4, -4, -70, 8, 96, -44, -22, -91, 93, 86, -128, 71, 21, -128, 127, -8, -87, 115, 57, -10, -128, 73, -37, -128, 120, 72, -117, 25, 6, -28, 46, -15, 127, -32, -128, 63, 117, -42, -29, 19, 44, 34, -106, -117, 127, 6, -115, 42, 124, -26, -128, 35, 13, -31, 34, 94, 34, -52, -75, 47, 98, -39, -123, 65, 119, -106, -62, 57, 42, 87, -120, -53, 127, -71, 17, 29, -20, -72, -110, 113, 59, -117, 108, 68, -122, -15, -20, 109, 73, -103, 2, -10, 49, 58, -128, 28, -45, -6, 41, 7, 72, -75, -9, -24, 88, -3, -128, 77, 78, -98, -39, 127, 1, -127, 31, 76, -1, 5, 27, -77, -53, -5, 109, -8, -127, -21, 127, -27, -29, 22, 24, 31, -45, 7, 11, 38, -30, 58, -79, -128, 127, 60, -128, -25, 127, -4, 43, -28, -128, 77, 52, -51, 69, -30, -54, 121, -58, -74, 127, -99, -44, 127, -65, -59, -23, -4, -56, 127, 9, -128, 49, -59, 127, 12, -88, 64, 52, -49, 3, 90, 17, -102, -107, 92, 20, 25, -19, 5, -15, -107, 127, -71, -128, 85, 27, -3, 36, 6, -54, 52, 61, -51, 27, -7, 0, -31, -126, 63, 72, 60, -41, -52, -38, 46, -3, -7, 66, -17, -7, 53, -88, -88, 127, -77, -5, 12, -36, 23, -14, 127, -125, -95, 86, 57, 80, -110, -115, -39, 111, 102, 14, -89, -95, -15, 115, 45, -29, 25, -122, 5, 47, -52, 105, -4, -81, 88, 11, -86, -76, 44, 12, -37, 95, 92, -128, -6, 127, -108, -47, 93, 38, -42, 10, -63, -52, 122, -15, -46, -75, 62, 100, -34, -128, 20, 127, -44, -82, -13, 64, -12, -8, 71, -22, -72, -24, 73, -85, -62, 127, 45, -128, 58, 8, 2, 127, -48, -34, -25, -56, -107, 47, 15, 20, 49, 30, 15, -128, -44, 127, 70, -63, -7, -7, -46, -77, -21, 0, 0, 64, 122, 39, -74, 17, -100, -26, 122, 45, -66, -82, 0, -14, 115, -27, 36, 2, -128, 58, 15, -4, 23, -58, -24, -15, 95, 79, -128, 71, 68, -107, -25, 44, -64, 95, 17, -128, 68, 108, 73, -8, -128, -72, -18, 127, 44, 15, -53, -53, 64, -29, -60, 56, 99, -128, 75, -4, -13, -29, -116, 64, 22, 6, 63, -6, -93, 89, 15, -36, 39, -55, -38, 64, 18, -59, 8, 108, -54, -38, 52, -20, 116, -18, -119, 28, 82, -92, 34, 65, -128, 105, 81, -99, -45, -37, 89, 2, 49, -90, 10, 77, -128, -28, 111, 62, -99, -34, -12, 41, 73, -4, 52, 26, -128, -22, 22, 68, 70, -128, -45, 113, 111, 28, -128, -80, -1, 99, 109, -128, 57, 110, -102, -88, 87, 2, -18, -14, -63, 127, 15, -128, 1, 76, 36, -22, 9, 91, -113, -104, 127, -18, 3, 106, -128, -96, -5, 23, 127, 59, -128, 52, -17, -2, -45, -111, 10, 93, 19, -55, 53, 43, -24, 43, -38, -128, 27, 127, 102, -92, -127, 68, 119, -128, -43, 127, -83, -56, 44, -76, 4, 111, -68, -2, 106, -128, 75, 68, -17, -105, 57, 24, -59, 68, -128, 103, 75, -128, 78, -5, -31, 127, -128, -93, 127, 5, -108, -31, -44, 95, 37, -42, 8, 8, -11, -110, 100, 12, -30, 77, -85, 22, 71, 42, 42, -49, -17, -30, -128, 28, 121, 18, -74, 34, -46, -63, 49, 2, 48, -1, -59, -59, -37, 108, 98, -94, 34, 0, -36, -3, 45, 62, 7, -41, -44, 91, -89, -52, 26, -29, -28, -30, 0, 55, 127, -54, -128, 14, 127, 26, 10, -105, -25, 127, -7, -83, -86, 32, 74, 22, 22, -38, -63, 71, -77, -98, 127, -8, 37, -72, 9, -1, -96, 2, 59, 49, -82, 80, 54, -95, -37, 68, -7, -70, 41, -4, 3, 102, 20, -81, -20, 45, 71, -91, -62, 0, 6, 27, 2, 38, -37, 10, 5, 48, 7, -126, 106, 105, -52, -36, 54, -100, 37, 39, -128, 77, -1, 63, -56, 30, 127, -87, -77, 49, 18, 1, 44, -128, -116, 53, 63, -3, 19, 102, -112, -128, 127, 127, -58, -39, -47, -2, 55, -49, 8, 74, 14, -128, -44, 127, 63, -78, -80, 26, -25, -56, 38, -7, -26, 71, 4, 29, 95, -128, -52, 127, -112, -73, 127, 58, -124, -100, 66, 86, 31, -120, 18, 49, -73, -32, 22, 0, 46, 91, -11, 19, 27, 14, 38, -128, -58, 44, 65, -6, -83, 48, -52, 4, 116, 71, -128, 37, -40, -58, 121, -42, 47, -94, 17, 127, -128, -128, 127, 93, -71, -9, -37, -3, 10, -25, -2, 98, 12, -91, -91, 125, 99, -128, -27, 71, -76, 36, 63, -106, -23, 127, 72, -128, -86, 96, 127, -73, -58, 98, 60, -103, -95, 34, 52, 61, 2, -108, 13, 20, -44, 107, -49, -87, -37, 80, 127, -120, -36, 9, -32, 123, -71, 48, 126, -128, -8, 72, -9, -77, -9, 60, -21, 40, 89, -128, -43, 94, -39, -70, 87, 103, -8, 34, 5, -18, -46, -13, -94, -115, 127, 21, -36, 119, -91, -56, -41, 57, 127, -95, 15, -45, 9, -15, 0, 93, -128, -7, -34, 18, 62, 46, -36, -95, 122, -27, -103, 46, 119, -51, -70, 80, 9, -74, -21, 119, 9, -69, 18, 23, -121, -2, 127, -128, -7, 127, -58, -115, -54, 107, 44, 6, -41, 47, -60, -104, 29, -9, 127, -83, -12, 49, 3, -8, -22, 13, -74, -5, 127, -100, 28, 13, -96, 127, -128, -70, 127, 0, -5, -96, -32, 41, 102, -81, -90, 51, -26, 87, 39, -92, 46, 15, -35, 43, 12, -64, 64, -66, -63, 127, -128, -37, 127, -31, -73, 86, -74, -103, 97, 74, -14, -128, -24, 93, -55, 34, 99, -51, -36, -47, 90, -38, -21, 47, 11, -14, -9, 70, -80, -38, 44, -5, -87, 43, -31, 36, 86, -99, -35, 0, -13, 108, 12, -42, 4, -1, 20, -82, -4, -53, 69, 41, -79, 40, 91, -35, -128, 127, 0, -45, 85, -128, -41, 127, 53, -80, 38, -47, 53, -44, -41, 71, -125, 20, -7, 79, -26, 23, -5, -63, 127, 13, 8, -83, -90, 108, 34, -65, 3, 76, -79, -128, 127, 57, -128, 48, -20, 58, -5, -128, 23, 111, 69, -103, -61, 68, 127, -98, -61, -37, 72, 48, -11, 75, -32, -71, -3, 44, -128, 9, 94, -55, 60, 35, -128, -66, 47, 36, -47, 14, 73, -29, -64, 127, 45, -128, 62, 13, -1, -46, -11, 63, 3, 7, -43, -22, 127, -54, -128, 5, 113, 82, -56, 20, -65, -4, 99, -57, 29, 40, -9, -93, 11, 127, -128, -82, 10, 76, 80, -35, 61, -93, -116, 72, 72, -13, 46, 8, -62, 69, 3, -107, 5, -46, 72, 86, -57, 12, -122, 17, 23, 26, 107, -128, -10, 127, -98, -2, 38, 22, -5, -121, 127, 19, -55, 42, -128, 36, 14, -6, 64, -7, 73, 22, -23, -15, -41, -36, -38, 37, -63, -4, 61, 7, 59, -128, -12, 127, 30, -128, 35, 26, -95, 121, 53, -114, -58, 108, 62, -47, -57, -21, -17, 18, 7, -28, -25, 127, 79, -65, -29, 55, -43, -128, 111, -19, -102, 54, 127, -77, -110, 127, -85, 20, 59, 17, -104, 6, 119, -39, -9, -122, -49, 127, 42, -44, -94, 61, 73, -11, 27, -128, 53, 127, -109, -65, 127, -31, -18, 77, -69, -96, 29, 80, -87, -90, 103, 0, -89, 43, -27, 58, 66, -83, 36, -73, 68, 83, -18, -17, -75, 11, 34, -23, -66, 121, 90, -128, -57, 112, -53, -115, -11, 127, 110, -105, -105, 29, 92, -48, 28, 96, -128, -49, 18, 39, 59, -110, -18, 47, 30, 52, 58, -128, 68, 18, -128, 127, 39, -62, 51, -3, 0, 28, -23, -34, -74, 66, -47, 28, 11, -12, 117, -128, -64, 106, 92, -53, 27, -89, -128, 64, 122, 53, -68, 0, 73, -44, -31, -31, -68, 20, -29, -56, 22, 109, 55, -54, -19, 51, -36, -5, 70, -105, -91, -26, 127, 127, -86, 36, -128, -2, 53, 2, 43, -12, 32, -70, -12, 3, -92, -108, 127, 22, -128, 17, 127, 68, -46, -39, -30, -42, -38, 11, 13, 14, -21, 22, -25, 127, 9, -128, 119, 64, -111, -25, 96, -75, -86, 56, 90, -31, -54, 85, -1, -40, 91, -20, -119, 51, 98, 0, -31, 57, 2, 12, -127, 25, 25, -128, 127, 0, -65, 34, 75, 1, 1, -19, -66, 96, 25, -128, -80, -21, 108, 62, -65, 7, 44, 32, -128, 0, 35, 22, 13, 47, 28, -107, 71, 18, -27, -15, 62, -66, -128, 127, 127, -128, -58, 104, -66, -60, 127, -2, -83, 46, 66, 28, 44, -42, -122, 98, 99, -92, -37, -35, 0, -43, 57, 26, -14, 23, 17, 44, -79, 73, -5, -128, 98, 81, -68, 25, 47, -98, -123, -28, 106, 89, -5, -7, -103, -82, 59, 127, 7, -128, -59, 127, -73, -4, 35, -47, 45, -128, 7, 125, 88, -3, -128, 40, 79, -41, 59, -49, -128, 95, 65, -29, 26, -86, -30, 81, -23, 25, 44, -8, 35, -21, 0, 2, 0, -128, 3, 14, -122, 127, 127, -128, -28, 127, 31, -128, -22, 98, -42, 29, -2, -122, 43, -11, -6, -27, 41, 127, -11, -71, -5, 62, -90, 0, 75, -121, 46, 35, -100, -42, 9, 39, -39, -25, 20, 2, -12, 127, 56, -23, 13, -96, -102, 26, 54, 35, -7, -60, 42, -17, 59, 29, -128, 17, -1, 96, 79, -128, -46, 127, -48, -39, 22, -82, 119, -5, -47, -57, -4, 10, 114, -35, -74, 10, -39, 127, -1, -14, -56, -109, 11, -27, 83, 23, -55, 117, -75, 29, 127, -128, 46, -47, -128, 37, 31, 127, -11, 14, -79, -128, 71, 4, -38, 127, -27, -41, 111, 13, -63, 23, 93, -100, 30, -23, -37, 6, -128, 125, -11, 25, 22, -128, -10, 53, 36, 18, -2, 68, 27, -113, 90, 48, -76, -106, 10, 87, 29, -73, -44, 6, -42, 21, 68, 127, -8, -123, -46, 94, -46, -47, 120, -55, -7, 63, -8, 59, -119, 31, 117, -88, -48, 23, -27, 31, 62, -21, -34, -90, 102, 65, -124, 55, 77, -27, 26, -81, -111, -13, -12, 3, 88, 61, -19, -83, -20, -21, 127, 44, -128, 68, 127, -51, -105, -23, 21, -35, -73, 127, 19, 24, 19, -62, 108, -90, -42, 104, -12, 32, -128, 21, 26, -51, 81, -23, 52, 12, -13, 24, -128, 34, 81, -128, -4, 127, -34, -23, 93, -79, -36, -36, -10, -52, 100, 53, -128, 90, -30, -100, 92, -12, 71, 75, -32, -9, -98, 60, 5, -103, 52, 72, -70, -82, 108, 104, -128, -66, 86, 104, 37, -128, -73, 28, -2, -10, 54, 48, 35, 17, -20, -73, 46, 39, 3, 46, -128, -46, 74, 4, 35, -64, -103, 127, -6, 3, 69, -110, -35, -28, 4, 127, -29, -69, -3, -25, 103, 1, 54, -24, -127, 38, 56, 105, -117, -80, 127, -122, 60, -2, -68, 89, -103, 54, 11, -59, 51, 47, 18, -27, 11, 55, -69, 25, -24, -66, -1, 46, 119, 40, -128, -128, 87, 77, 96, -36, -128, 65, 75, -128, 74, 4, -87, 127, 10, -38, -103, 106, -1, -78, 71, 18, -28, 7, 38, -47, -64, 38, 29, -128, 90, 51, -128, 127, 127, -128, -49, 10, 25, 127, -128, -93, 127, -4, -128, 8, 127, -54, -76, -32, 63, 127, -21, -124, -1, 23, -18, 121, -128, 21, 127, -83, -124, 77, 81, -128, 116, -15, -128, 127, 120, -81, -128, 117, 105, -100, -64, 73, 40, 0, 34, -54, -9, 14, 13, -18, -128, 43, 68, -116, 62, 21, -4, 117, -92, -107, 127, -23, -113, -9, 123, 4, -124, 127, 112, -128, -90, 54, 49, 127, -128, -56, 80, 40, -47, -85, 32, -35, 108, 57, -115, -25, 80, 100, -128, 31, 21, -128, 19, 65, -25, 103, 64, -122, 102, -10, -64, -37, 48, 21, -125, 107, 106, -48, -10, -87, -128, 127, 23, -21, 40, -53, -19, -61, 54, 30, -69, 47, 49, -56, -81, 69, 35, -14, -20, -45, -15, 72, 61, 29, -102, -23, 127, -128, -24, 123, -112, 35, 68, -45, 41, -73, -88, 127, 8, -35, 15, -20, 39, -117, -65, 116, 97, -36, -56, -70, -76, 85, 127, -21, -42, -104, 0, 87, -87, -64, 127, -15, -36, 54, -15, 0, -56, 122, -58, 1, 75, -39, 18, -106, 39, 127, -128, -4, 102, -83, 70, 18, -128, 73, 2, -41, 115, 0, -128, 29, 127, -128, -128, 124, 45, 5, 78, 21, -35, -128, 64, 42, -128, 51, 127, -122, -39, 127, -128, -117, 110, 91, 46, -53, 6, -99, -49, 90, 59, -12, -71, 32, 11, -19, -38, -87, 24, 42, -54, -41, 113, -29, -26, 127, 9, -51, -128, 14, 100, -112, 80, 13, -128, 127, 119, -7, 27, -90, -66, 127, -103, -128, 127, 68, 39, -128, 29, 54, -89, -30, 19, 17, -54, -8, 123, 127, -108, 25, -37, -5, 127, -128, -128, 127, 124, -59, 0, 2, -110, -60, 103, -53, -1, 2, 63, 26, -128, 91, 49, -35, 54, -122, -12, 127, -128, -43, 127, -20, -26, -86, 21, 72, -80, 34, 43, -102, 13, 51, -128, 65, 127, -69, 47, -60, -21, 100, -31, -119, 8, 24, 41, 18, -91, 65, -28, 0, 10, -77, 27, -51, 37, 9, -5, 127, 31, -121, -107, 53, 85, -51, -73, 40, 114, -73, -13, 125, -128, -35, 127, -2, -17, 47, -128, -64, 77, 37, -104, 62, 127, -125, 46, -14, -75, 69, -57, -31, 106, -18, 18, -5, -25, -64, 40, 82, -128, 62, -18, -59, 17, -37, -15, 5, -17, 10, 91, 20, 42, 13, -79, 41, -70, -26, -4, 55, -2, -52, 21, 68, 127, -128, -79, 127, -35, -39, -11, 66, -25, -19, 5, -40, 127, -55, -35, 102, -15, -107, -23, 32, 64, 46, 29, 26, -128, -121, 88, 11, -26, 103, -74, -60, 127, -11, 63, -93, -7, 41, -20, -35, -9, 127, -85, -38, -36, -77, 31, 111, -35, -30, 127, 57, -128, 21, 86, -97, -102, -43, 114, 15, 18, 35, -15, -6, -123, 54, 57, 14, 94, -128, 19, 111, -128, -17, 41, -49, 54, 34, 54, 46, -128, 45, 107, -115, 65, -24, -12, 105, -74, -55, -27, -11, -52, 119, 127, -128, 13, 36, -123, 72, 73, -105, -32, 96, 23, -31, 44, 68, 27, -58, -72, 97, -23, -128, 31, 6, 22, 12, -66, -41, 115, 55, -98, 95, 14, -128, 127, -18, -113, 23, 21, 127, -128, 23, 44, -61, -18, 92, 37, -128, 40, 127, -121, 27, 5, -81, 31, -3, 120, -82, -9, 38, -26, 113, -99, -4, 127, -128, 23, 52, -128, 43, 127, -70, -128, 29, 60, 36, -107, 109, 41, -73, 74, -34, -51, 48, 66, -28, -108, 2, 82, 22, 35, -97, -51, 127, -113, -58, 22, -121, 127, 6, -78, 127, -56, -22, 113, 1, 2, 34, -51, -105, 5, -7, 19, 127, -128, -54, 110, -71, -58, 13, -37, 127, 61, -91, 104, -7, -128, 95, 55, -11, -56, -128, 123, 42, -8, 40, -102, 38, 38, 43, -72, -128, 41, 127, -41, -103, 86, 37, 12, -15, 44, 1, -42, -42, -44, 29, 107, -17, -71, 21, -22, 26, 36, -96, -71, 32, 102, -26, 64, -11, -128, 127, -6, -127, 127, -45, -8, -12, 39, -6, -22, 78, 2, -68, 3, 127, -47, -46, -25, -75, -55, 113, 102, -60, 13, 20, 3, -85, 37, 59, -95, -94, 25, 94, -38, -64, 59, 127, -88, -59, -22, -66, -11, 127, 10, -9, 86, 2, -27, -124, -61, 73, 127, 35, -128, 0, 94, -128, -74, 105, 82, -23, 3, -45, -112, 127, 31, -55, 98, -11, -121, 43, 105, -128, 26, -32, -113, 120, -58, 19, 127, -126, -60, 93, 100, -26, -99, 15, 26, 4, -76, -30, -11, 86, 69, -126, 56, 102, 35, -44, -55, -45, 5, 18, 9, -7, -42, 85, 63, -69, -53, 21, -3, 65, -81, -45, 44, -22, 115, 65, -128, -105, 39, -28, 127, 63, -124, 24, 21, -82, 127, 111, -128, -8, -54, 72, 124, -103, -1, 37, -128, -47, 26, 64, -26, -42, 17, -18, 127, -61, -128, 127, -21, -128, 127, 103, -79, 54, -73, -18, -1, -117, 105, 21, 18, 44, -64, -7, -17, -59, 2, 12, 42, -10, 76, 8, -59, 83, 21, -100, 23, 110, -128, 45, 4, -128, 127, 117, -128, -97, 111, 0, -27, -18, 71, -20, 31, 0, -21, 11, -90, 127, -22, -17, -3, -91, -6, 127, -53, 25, 26, -22, 127, -128, 20, 98, -105, -20, 36, -59, 26, 107, -64, 25, -74, -128, 12, 116, 10, -47, 122, -52, -41, -45, -62, 113, 7, -71, 49, 0, -57, 83, -24, 40, 127, -14, -19, -115, 8, -18, 21, 28, -94, 4, 23, -5, 14, -3, 107, 15, -20, 28, 8, -72, -10, -55, 8, 127, -128, -95, -3, 1, 127, -35, -115, 123, -44, 23, 127, -42, -128, -8, 127, -103, -6, 10, -64, -2, 12, 36, 15, 23, -117, 36, 109, 17, -26, -35, 13, 30, 10, 4, -121, -43, 127, -57, -116, -27, 9, 4, 92, 5, -6, 79, -52, -20, 57, 65, -31, -87, -43, -9, 91, 21, -128, 59, 41, -5, 17, -127, 74, -3, 39, 98, -53, 46, -128, 26, 127, -128, -122, 68, 59, 49, -47, -128, 70, 11, -61, 9, 87, 39, -2, -12, 64, 42, -128, -35, 43, 20, -12, 74, 49, -128, 26, 2, 65, 69, -128, 45, 122, -105, -77, 2, 127, 15, -128, 18, 32, -15, -14, 119, 11, 9, -56, -69, 59, -53, 45, 58, 0, -128, -12, 55, -107, 127, 52, -128, 45, 81, 34, -61, -12, 127, -70, -25, -32, -10, 127, -43, 3, -38, -74, 60, -64, 70, -52, 3, 9, 0, 61, -21, 54, 41, -128, -7, 127, -128, 20, 2, -15, 43, -56, 1, -8, -77, -55, 116, 94, -112, -68, 104, 2, 45, -70, -13, 106, -115, -17, 119, -83, -128, 127, -23, -128, 127, 127, -128, -128, 127, 65, -128, 39, 14, 24, -8, -90, 127, 96, -128, -107, 35, 105, 78, -113, -106, 70, 127, -38, -128, 85, 70, -98, -3, 52, -9, -62, 24, 52, -34, 6, -65, 25, -1, -40, 46, -46, 92, 3, -128, 127, 37, -98, 85, -68, -15, 121, -3, -26, -66, -98, 26, 127, -12, -128, 34, 127, -52, -128, 42, 110, 15, -25, -60, 58, -75, -6, 5, 22, -9, -116, 127, -8, 10, 1, -32, 22, -65, 11, -36, 27, 59, -11, -2, 48, 36, -128, 76, -12, -106, 75, 103, -58, -128, 90, -35, -12, 38, -18, 6, -3, 53, 112, 18, -97, -32, -7, 82, 45, -2, -111, -71, 58, 69, -79, -72, 111, -52, -34, 71, 25, 34, -18, -25, 79, 23, -29, -95, -82, -41, 69, 58, 4, 23, -68, -86, 127, 107, -128, 49, 106, -119, -27, -13, -39, 49, 63, 30, -8, 57, -59, -128, 98, 75, 26, -18, -41, 3, 44, 20, -44, -44, -65, -32, 127, 10, -122, 91, 121, -104, -55, 46, -25, 62, -10, -29, -83, 59, 127, -103, -37, -66, 2, 10, 18, 23, 0, -28, 32, 38, -1, -12, -37, 115, -56, -53, -61, 52, 29, -128, 127, 116, -116, -30, -5, 68, 79, -95, -25, 72, 35, -112, 15, 31, -94, 28, 61, -100, 6, 89, -56, -1, 78, -61, -69, 32, 38, 53, -107, -114, 127, -7, 11, 6, -37, 37, -108, 52, 96, 49, -71, -12, -22, -48, -8, 44, 127, 8, -23, -25, -51, -40, -20, 0, 60, 55, 26, -59, -37, -78, 21, 48, -75, 30, 23, 75, 20, -52, -34, -28, 0, 91, -87, -11, 36, -93, 63, -21, -36, 8, 114, 57, -36, -64, -87, 29, 127, 85, -30, -83, 49, -20, -29, -30, 11, 26, -128, 42, 127, -28, 6, -21, -121, 115, 107, -90, -128, -11, 83, -27, -4, 6, 37, 127, -106, -19, 9, -107, 110, -58, 8, 116, -68, -27, 91, -61, 5, -54, -11, 127, -76, -6, 73, 23, -92, 38, -64, -26, -11, -8, 127, -65, 29, 7, -73, -30, -42, 94, 48, -128, 85, 47, -43, 9, 26, 40, -44, 26, -11, -26, -29, -44, -31, 54, -52, 76, 48, -107, 43, 38, -83, -10, 20, -85, 127, 92, -123, -37, 3, 119, -24, -104, -12, 124, 86, -128, 22, 41, 39, -32, 25, 3, -71, -7, 22, 97, -127, -108, 127, 61, -109, 100, 39, -60, -128, 53, 38, -111, 127, 36, -128, -45, 124, 19, -115, 29, 32, 48, 65, -85, -128, 97, 77, -56, 82, -54, -128, 127, 17, -128, 25, 127, -57, -113, 87, -46, 89, 81, -126, 93, -70, -38, 1, 25, 127, -124, -102, 47, -30, -68, 125, -14, 28, 6, -27, 100, -45, -128, 27, 127, -104, -128, 126, 29, -69, -20, 31, 10, 63, -62, -79, 3, 56, 68, 27, 23, -15, -40, -128, 127, 32, -28, -21, -89, 17, -42, -13, 127, -31, 10, 106, -95, -96, 10, 127, -22, -10, -28, 31, 41, -86, -53, 52, -36, 20, 74, -4, 1, -1, 65, -45, -110, 43, 91, -48, 20, 41, -31, -44, 49, 5, -123, -34, 69, 37, 55, 77, -128, -120, 115, 64, -59, 59, -78, -51, 69, -1, -24, -116, 44, 9, -1, 80, 46, -68, -114, 73, 127, 37, -128, 37, 45, -94, -37, 82, 127, -128, 18, 31, -105, 93, 64, 57, -46, -128, 49, -9, 0, 127, -128, -128, 127, 48, -72, 42, -15, 30, -85, -28, 71, -55, -31, 89, 32, -80, 17, 9, -27, -8, 12, 51, 75, -79, -37, 29, -44, -30, 26, -7, -81, 93, 24, -90, 1, -41, 110, 127, -17, -128, -44, 59, -32, 110, -86, 47, 19, -61, 52, -5, -38, -122, 93, 1, 0, 14, 3, 127, -25, -125, -53, 89, 114, -72, 34, -85, -70, 127, 51, -93, 8, 0, -31, 10, -113, 121, 9, -83, 52, 68, -92, -17, 127, -47, 19, -66, 7, 49, -112, -7, 83, -20, 78, 2, -48, 103, -79, -87, 53, -21, 14, 17, -9, -18, -2, 63, 57, 1, 6, -47, -117, 127, -75, -128, 107, 97, -45, -77, -30, 38, 60, 8, 54, -60, 52, 31, -128, -18, 104, 57, -45, -39, -70, -49, 99, 73, 6, -1, -71, 21, 106, 0, -63, 36, 54, -128, -6, 14, -75, 111, 8, 15, -41, -87, 0, -21, 108, 3, -41, 18, 68, 95, -64, -7, 73, -128, -80, 87, 25, 30, -88, -9, 32, 41, 18, -96, -66, -19, 81, 6, 46, 123, -128, -128, 42, 18, -11, 109, 14, -25, -32, -61, 71, 93, -76, -35, -27, 38, 6, 7, 63, -73, -8, 103, -39, 15, 0, -100, -4, 45, 127, -128, -10, 127, -128, 28, 6, -119, 127, 27, -128, 62, 127, -87, -2, -72, -115, 127, 111, -113, -18, -8, 3, 127, -128, 12, 127, -128, -93, 127, -55, -128, 13, 127, -8, -126, 127, -37, -18, 49, -2, 51, -88, 6, -27, 68, 79, -128, 41, 3, -29, -20, -32, 127, 89, -128, 15, 64, -45, -82, 8, 98, -91, 20, 35, -97, 116, -46, -87, 87, 4, -53, -82, 116, 94, -117, 28, -13, -32, 26, -38, 124, -41, -35, 89, 48, 39, -95, -27, -3, 13, -21, -122, 124, 127, -92, -127, 73, 53, -30, -69, 66, 94, -128, 29, 1, -45, 14, -39, 109, -5, -42, 32, -7, -49, -60, 52, 127, 26, -128, 0, 47, -39, 60, -20, -78, 127, -6, -6, 21, 1, -47, -94, 103, -13, -104, 77, 127, -128, 72, 37, -98, 24, 39, 80, -74, 9, -27, -76, 43, -42, 73, 46, -45, -61, 28, 93, -96, -120, 89, 121, -128, 51, 20, -53, 29, -77, 21, 123, 6, -102, -18, 99, 102, -128, 36, 68, -128, -19, 127, 27, -68, 70, -74, -73, 9, -35, -6, 75, -8, 79, 0, -127, 124, -9, 6, 106, -55, -128, 82, -46, -42, 57, -126, 70, 39, 60, 94, -90, -122, 104, -59, 5, 127, -123, -69, 108, 24, -82, -12, 60, -13, -10, -34, -77, 23, -21, 0, 126, 32, -128, 90, 127, -128, 0, 43, -59, 88, -48, -105, -26, 22, 30, -23, -64, 108, 47, 39, -62, 9, 15, 4, -9, 11, -37, -80, 34, -90, 108, 115, -63, -10, 43, -38, -106, 11, 127, 18, -96, -26, -79, 34, 127, -88, 4, 108, -128, -92, 127, -12, -89, -13, -2, 97, -46, -28, 13, -44, 69, 77, 64, 31, -96, -38, -3, -8, -31, -19, 20, 29, 98, -65, -89, 56, 75, -90, -53, 127, 0, -128, 127, 91, -128, -28, 4, -8, 87, -21, -55, 127, 83, -128, 31, -8, 3, -11, -45, 127, -80, 5, 28, -127, -53, 97, 78, -17, 0, 57, -83, 1, 127, -128, -87, 127, -41, -83, -21, 52, 74, -88, 43, -28, -7, 27, -28, -9, 18, -39, -71, 127, 112, -82, 4, 85, -128, -60, 70, 46, -46, -7, 85, -128, 72, -10, -128, 41, 61, -7, 92, -59, -52, 125, -81, -61, 122, 72, -78, -51, 35, 68, -113, 2, 24, -102, 60, 35, 21, -62, -96, 127, 71, -18, -113, -39, 127, -104, 0, 31, -66, 81, -24, -82, -14, 89, 34, -89, 20, -41, 55, 11, 31, -25, -128, 68, 29, 40, 62, 49, -30, -6, 59, -110, 13, -52, -128, 127, 1, 47, -48, -15, 119, -71, -66, -80, 28, 125, -19, 4, 114, -127, -128, 127, 1, -110, -7, 38, 127, -128, -52, 119, 38, 1, -128, 62, 103, -126, 19, -36, -72, 127, 93, 39, -99, -120, -32, 86, 127, -58, -62, 81, 6, -11, 39, -128, -77, -3, 102, 25, -128, 43, 127, -70, -128, 25, -38, 122, 49, -57, 79, 4, -91, 26, 51, -32, 52, 10, -105, 53, -6, -128, 127, 6, -128, 127, 31, -99, 127, -61, -28, -2, -11, 116, -104, 31, 94, -110, -3, -43, 65, 26, -32, 6, -128, 27, 127, 106, -128, -119, 127, -9, -96, 77, 1, -42, -2, 39, 79, -93, 25, 40, -93, 49, -69, 41, 32, 35, -71, -2, 127, -14, -128, -3, -5, -73, 17, -56, 43, 12, 12, -20, 13, 100, 11, 12, 47, 36, -110, -21, -15, -77, -8, 53, 117, -83, -59, -32, 127, 11, -42, 127, -128, -128, 127, 3, -55, 106, -54, -18, 113, -51, -11, -35, -100, 40, -20, -42, 48, 32, 86, -6, -46, 65, 78, -128, 25, 9, -128, 127, 23, -128, 110, 66, -112, 9, 77, 48, -86, -123, 75, -7, 25, 21, -71, 113, 18, -93, 64, 56, -32, -11, -99, -39, 60, -52, 30, 46, -74, 99, -23, -6, -36, -95, 70, 5, 96, -48, -87, 18, -12, 127, 3, -128, -27, 127, 114, -14, -123, 29, 80, -128, -8, 127, -5, -128, -54, 31, 60, 20, 87, 68, -128, -128, 127, 66, -128, 73, 24, -31, 42, 43, -57, -128, 95, 94, -128, 68, 80, -128, 95, -59, -46, 42, 52, 127, -128, 35, -32, -49, 82, -128, 28, 92, -75, -32, 127, 12, -128, 44, 20, -110, 60, 122, -63, -36, 32, -34, -11, 81, 56, -128, 32, 127, -117, -69, 127, -34, -82, 113, -91, 6, -22, -55, 96, -128, 127, 23, -72, -27, 36, 127, -128, -57, 71, -15, 52, 59, -17, -122, -4, 40, -79, 26, 12, -1, 127, -85, 7, 86, -128, -34, 60, -19, 59, 113, -117, 0, 127, -9, -37, 20, -26, -128, -28, 11, 38, -21, 81, 13, -128, 75, 24, -29, 57, 30, 0, -2, -9, 2, 51, 13, -37, -83, 38, 14, -6, 127, -128, -4, 127, -28, 14, -109, 24, 126, -99, -128, 127, -28, -111, 9, 14, 96, -29, -81, -55, 127, 56, -71, 9, -40, -12, -63, 75, -18, -41, 105, -100, 11, 51, 40, 14, -122, -24, 46, -22, 32, 103, -103, 14, 127, -104, -124, 86, 62, -64, 27, 32, 30, -15, -128, 0, 127, -54, 35, 105, -64, -59, 47, -62, -1, 86, -79, 64, 17, -38, 69, -108, -120, 127, 87, -128, -125, 127, 88, -68, -65, -32, 7, -65, 112, 12, -66, 45, -1, 0, -71, 127, 81, -28, -87, -65, 59, 25, -7, -107, 35, 29, -57, 104, -42, 39, 127, -128, 42, 44, -10, -66, -15, 127, -128, -57, 9, -13, 127, -30, -19, 90, -59, -83, 66, 7, 34, -70, -108, 32, -19, 77, 18, -41, -18, 20, -8, 94, 26, 23, -13, -128, 127, 127, -128, -128, 96, -22, 39, -3, -4, 12, 55, 120, -80, -35, -18, -39, 52, 22, -45, 30, 93, -39, 22, -125, 24, 3, -28, 82, -128, -37, 105, -7, -107, 120, 2, -49, 96, 30, -21, -109, 90, 22, 15, 3, -6, -7, -29, 39, 15, -44, -113, 116, 112, -128, 1, 127, -128, 8, -6, -85, 116, 57, -100, 41, -22, -53, -13, 41, 127, -85, -30, 55, -21, 12, -125, -18, 127, 28, -128, -3, 127, -105, -78, 104, -10, -82, 13, 97, -123, 17, 6, 0, 68, -87, 39, 12, 43, 14, -104, 59, -27, -128, 88, 112, 29, -42, -63, 42, -10, -42, 36, -56, 86, -53, -128, 86, 17, 70, -49, -56, 76, -37, -58, 113, 58, -28, -31, -42, -10, 60, -23, -66, 115, 54, -113, 0, 12, 18, -1, 12, -30, 36, -7, -128, 127, 1, -82, 9, 78, 45, -53, -36, 10, 105, -125, -71, 82, 1, 30, 64, -95, -128, 42, -10, 73, 74, -15, -71, -51, -11, 99, 66, -14, 85, -71, 6, -63, -114, 23, -11, 95, 115, -56, -47, 32, 49, -128, -68, 95, -92, -29, 127, -86, -27, 127, 13, -111, -54, 127, -21, -72, 82, -104, -42, 127, 20, -42, -111, -82, 127, 22, 9, 57, 6, -10, -92, 63, 52, -128, -58, 127, -8, -128, 113, -8, -128, 127, 34, -32, 45, 56, -73, -93, 127, 61, -128, 28, 24, -115, 127, -70, -44, 127, -8, -5, -65, -56, 62, -41, -56, 127, 69, -32, -128, 0, 127, -121, -54, 4, 42, 127, 17, 0, -120, 20, 63, -86, 47, -128, 36, 127, -128, 26, 39, 35, -26, -15, -23, 4, 125, -90, 0, 48, -122, 63, 7, 1, 127, -94, 37, 11, -108, 98, -23, -30, 113, -128, -69, 125, -78, -34, 35, -35, -51, 46, 127, -88, -123, -22, 112, 127, -120, -40, 4, -6, -24, 18, 29, -119, 127, 18, -100, 86, -69, -79, 61, 15, -60, 127, 97, -107, -48, -49, 53, 40, -4, 45, -41, 51, 10, -81, 11, 87, 18, 9, -77, -128, 35, 106, -82, -32, 127, 0, 8, 59, -52, -88, -112, 122, 5, -3, 10, -75, 127, 14, -2, -32, -88, 0, -12, 80, 100, -128, 22, 127, -128, -82, 127, 3, -17, 81, -2, -43, -68, 46, 17, -110, -73, 106, -32, -56, 99, -57, 89, 32, -128, 93, 127, -88, -103, -5, 38, -37, -3, 21, 94, -1, -68, 70, 41, -57, -36, 83, -98, -94, 103, 80, -58, 27, -8, -51, 2, -128, 127, 43, -95, -22, -46, 69, 48, 0, 23, 80, -10, -128, -44, 91, 9, 71, -35, -93, 53, -65, -36, 117, -14, 63, 3, -29, 81, -3, -44, -128, 99, 35, -87, 3, -18, 53, 23, 61, -109, -97, 127, 34, -56, -88, -54, 127, 124, -97, -96, -4, 32, 11, 68, 48, -86, -78, 59, -2, -71, -17, 56, -14, 28, -38, -5, 4, 21, 15, 34, 95, -92, 24, -15, -128, 95, 74, 0, 62, -128, -51, 25, 19, 127, -103, -73, 60, 14, -53, 30, 127, -77, -105, 119, 127, -128, -78, 127, 52, -73, 15, -1, -121, 9, 127, -79, -89, 68, -34, -59, 58, 63, -77, 114, 7, -128, 35, 36, 62, -28, -87, 6, 85, -11, -65, 36, 30, 35, -18, -63, 6, -32, 96, 30, -24, 43, -42, 68, 68, -82, 40, -73, 20, -9, -128, 38, 11, 41, 36, 73, 0, -23, -77, -97, 127, -1, -62, -1, 38, 102, -109, 42, 57, 13, -88, -112, 60, 60, -49, -55, 25, -44, 71, 5, -81, 116, 1, -72, 127, 63, -128, 2, 45, -86, 93, -27, -39, 19, -23, -2, 85, 89, -128, 1, 109, -90, 39, 127, -36, 21, -126, 34, -34, -47, 34, -110, 65, -1, 43, -20, 73, 60, -23, -76, 18, 58, -97, -22, 45, 61, -36, -21, -31, 0, 126, 32, -59, 2, 12, -49, -11, 87, -59, -35, 37, -58, 41, 55, -26, -76, -111, 52, 127, 9, -30, 2, -77, -123, 127, 114, -65, -52, -91, 93, 127, -128, -14, 70, 32, -8, -128, 70, 41, -23, -8, 86, -49, -128, 127, 80, -82, 34, -24, -90, 83, -48, -114, 127, -26, 21, 87, -47, -40, -2, 80, -128, 75, 15, -58, 107, -28, 3, -60, 61, -30, -63, 127, -116, 10, 58, 8, -42, -91, -5, 25, 127, -99, -53, 110, -86, -3, 13, -125, 113, 127, -89, 9, 37, -32, -20, -43, -12, -53, 96, 3, -78, 68, -76, 43, 30, -7, 45, -8, -66, -128, 64, 39, -47, -27, 123, 49, -38, -58, -35, 103, -83, -75, 77, 127, -114, -123, 116, 25, 7, 17, -116, -26, 49, 7, -26, 87, 31, -128, 89, 119, -126, -76, 127, 5, -111, 96, 95, -122, -128, 70, 127, -82, -10, 62, -116, 70, 80, -5, -62, -57, 17, -20, 65, 26, -18, 65, -43, -128, 127, 0, -82, 127, -87, -66, 10, 31, 23, -111, 111, 19, -43, 54, -22, -22, -110, 98, -1, -18, 87, -57, -77, 72, 105, -21, -58, -58, 49, 52, -48, -10, -93, -88, 127, -20, 28, -36, -128, 54, 47, -63, 85, -1, -3, 60, -60, 112, -79, -13, 85, 8, -40, -128, 126, 66, -128, 78, -22, 54, 85, -61, 37, -5, -113, -34, 127, 56, -77, -110, -72, 127, -31, 9, -30, 8, 60, -86, 114, -15, -68, 15, 2, 44, 19, -63, -71, 57, -34, -83, 107, 53, -114, -38, 58, -74, 114, -2, 30, 26, -111, -5, -31, 94, -43, -52, 99, -19, 83, 14, -128, 59, -4, 20, 60, 24, -48, -4, 77, -81, -57, 0, -17, -12, 111, -2, -51, 24, 38, -26, 20, 111, -43, -128, 22, 104, -34, -111, 127, 38, -90, -51, 66, 88, -41, -26, -74, 127, -79, 12, 56, -128, 11, 7, 43, 79, -1, 18, -58, -112, 31, -31, -27, 127, -51, -8, 63, -83, 102, -40, 3, 0, -87, 63, 91, -96, -128, 65, 10, -30, 39, 40, 25, 2, 80, -94, -68, 124, -106, 36, 127, -80, -128, -17, 73, -8, -65, 109, 91, 24, -90, -49, 27, 14, 10, -98, 120, 1, -34, -64, 14, -5, -17, 34, 2, 57, -58, -28, -44, 70, -2, -68, 0, 2, 64, 32, -12, 25, -19, -66, 57, 46, 27, 79, -95, -111, 25, -7, 53, 127, -75, -124, 127, 87, -99, -12, -39, 38, 98, -87, -82, 102, 24, -89, -88, 95, 124, -111, -31, -79, 18, 127, -38, -108, 63, 58, -35, -128, 98, 7, -1, 17, -114, 127, -122, 23, 111, -128, 98, -14, -7, 4, -91, 27, 70, 3, -73, 54, -100, 53, 120, -89, 61, -68, -128, 93, 127, -42, -52, 55, 4, -25, -114, -60, 111, -39, -38, 1, 42, 11, -2, 32, -13, 89, 49, -103, -52, -17, 105, 30, -128, 45, 127, 51, -66, 15, -17, -63, 12, -66, 2, -9, 69, 32, -72, -10, 0, 72, -53, 41, 73, -28, -88, -88, 65, 121, -43, 6, -55, -85, 43, -56, 127, -15, -128, 122, -35, 32, 12, -11, -36, -14, 127, 22, -128, -57, 13, 56, -28, -28, 91, 49, -64, 5, -5, -128, 127, 104, 7, -114, -122, 53, 25, -18, 9, 61, 55, 10, -106, 112, -10, -128, 127, -32, -107, 127, 55, -95, 7, 66, -97, -85, 124, 35, -120, 86, 74, -128, 48, 88, -128, 76, 102, -114, 51, 102, -24, -56, -36, -87, 23, 111, -39, -77, 83, 71, -128, -1, -22, 73, 20, -108, -13, 112, 109, -128, 43, -4, -91, 48, 52, -7, -71, -29, 107, -29, -107, 92, 70, 2, 0, -63, -31, -38, 54, 10, 5, 112, -39, 13, 22, -128, -88, 127, 127, -128, -121, 127, -25, -28, 34, -115, -30, 121, 4, 35, 83, -75, -35, 3, -27, -68, 103, 83, -112, 0, -54, -61, 76, 102, -49, -119, 127, 40, -128, 87, 56, -86, 34, 79, -121, 37, 127, -128, 0, 1, -83, 52, 89, 26, 49, -98, -128, 127, 127, -110, -71, 95, 6, -1, 1, -3, -92, -47, 42, -43, -1, 73, 54, 25, -43, -25, 94, -123, 48, 45, -111, -40, 105, -28, -6, 127, -128, 27, 112, -128, -37, 8, 89, 114, 0, -68, -34, -85, 41, 127, -128, -113, 43, 115, 53, -6, -64, -40, 105, -63, 15, -11, -98, 114, -38, -69, 41, 31, -47, -63, 64, 56, -60, -4, 25, -52, 85, 127, -128, -26, 109, -87, 38, -43, -114, 98, 104, 4, -128, 63, -18, -115, 19, 82, -44, -7, 6, 2, 22, -71, 127, 38, 17, -95, -112, 44, 42, -28, -35, 98, 86, 66, -128, -20, 24, -69, 72, -49, -57, 127, -30, -65, 7, -4, 15, -69, 127, -21, -68, 127, -65, -104, 79, -42, -41, 117, -37, 0, 77, -45, -63, 18, 23, -13, -45, 59, -86, -6, 127, -128, -68, 127, -35, -66, -27, -17, 86, -91, 5, 48, -126, 127, 87, -52, -60, -100, 71, 55, 82, -46, -128, 62, -64, 88, 3, -99, 127, -79, -70, 113, -32, 44, 47, -19, -31, 26, -38, 22, 119, -39, -125, 37, 90, -31, -21, 31, -100, -128, 127, -49, -22, 127, -31, -52, 42, -25, 70, -55, -57, -5, 26, 93, 28, -83, -75, 40, -92, 86, 18, 37, 39, -105, 107, -57, -92, 91, -53, -30, 103, 38, -48, -78, 4, 111, 48, -128, -56, 126, -46, 31, 113, -128, -19, 127, -70, -97, -30, 37, 127, -18, -79, -18, 111, -21, -65, 17, 37, 63, -23, -18, -42, -65, 61, 107, 42, -86, 1, -23, 42, -12, -128, 127, -37, -6, 81, -97, 79, 2, -23, 11, -10, 76, -14, -57, -91, -75, 117, 91, -15, -59, -110, 127, 14, -54, 87, -91, -95, 52, 86, -92, 11, 98, 26, 5, -71, -40, -46, -23, 124, 75, -15, -44, 1, 11, -128, 72, 82, -22, 9, -117, 109, 79, -128, -17, 30, 69, 37, -66, -70, 127, 20, -69, 69, -98, -56, 127, 6, -110, -24, -14, -28, 116, 86, -28, -68, -4, 31, 21, -29, 6, 126, -122, -55, -43, 19, 121, 19, -96, -128, 127, -15, -103, 112, 20, -17, 44, 19, -128, -58, 127, -25, -90, 74, 103, -128, 12, 91, -91, 28, 63, -53, -27, -46, 47, 74, -32, 13, -89, 61, 63, -128, 94, -48, -21, 109, -64, 58, -92, -21, 127, 15, -15, -107, -55, 89, -45, -43, -36, 63, 127, 20, -128, -85, 127, 45, -15, -21, -89, -61, 7, 127, -18, -94, -56, -34, 127, 62, -128, -69, 81, -24, -42, 38, 30, 52, 87, -15, -1, 78, -115, -20, 102, -68, -112, 88, 22, -123, 38, 91, 0, -128, 45, 127, -96, -15, -14, -73, 52, -28, 6, 94, -55, -42, 122, 1, -128, 59, 24, -128, 111, 68, 14, 15, -128, -52, 73, 36, 8, -83, -12, 9, -36, 30, -29, 66, 127, -89, 28, 11, -78, 68, -120, 99, 14, -128, 112, 21, 34, 93, -93, -18, 11, -32, -32, 28, 60, 32, -89, -114, 127, 44, -128, 106, 64, -128, 14, 37, -2, -3, 59, -82, 31, 124, 10, -128, -7, 113, -125, 61, -19, 19, -4, 2, -20, -31, 25, 45, -1, -98, 127, -94, -5, 2, 18, 52, -128, 30, 58, 42, 20, -77, 0, 80, -128, 21, 85, 42, -99, 8, 93, -113, 21, 94, -115, 7, 55, -83, 48, 56, -128, -14, 127, -9, -19, 23, -108, -114, 22, 109, 112, -128, -110, 119, 80, -62, -56, 24, -17, 39, -10, 81, -40, -128, 127, 35, -128, 21, 127, 61, -117, -128, 90, 8, 40, 63, -128, -55, 108, 20, 52, 24, -92, -29, -40, 0, 65, 52, -18, 82, -108, 13, 127, -128, -122, 116, 83, -109, -59, 90, -40, -18, 95, 5, 22, -22, -113, 71, 62, -10, -65, -29, 18, 0, 89, -65, 36, -45, 29, 10, 1, 127, -128, 14, 0, -102, 91, 56, -26, 25, -49, -22, -3, 51, -23, 24, 22, -128, 89, 92, -128, 29, 56, -124, 28, 109, 30, -128, -77, 68, 29, 112, -21, -97, 121, -57, 22, 11, -128, 40, 4, -34, 127, -4, -128, -5, 26, 35, 45, -75, -51, 93, 100, -39, 0, -32, -75, 38, -10, -3, 62, 49, -54, -108, -2, 30, 35, -20, 14, 76, -23, 13, 70, -23, -128, -64, 127, 36, -30, -17, -31, 96, 64, -89, -89, 71, 30, 22, -125, 68, 8, -55, 117, -76, 23, 65, -9, -128, 90, -5, -57, 59, 10, 47, -128, 76, 125, -62, -40, -90, 111, 106, -128, 34, 18, -81, 61, 60, -65, -56, 123, -55, -76, 18, 64, 127, -112, -90, 30, -53, 66, 119, 0, -75, -20, 43, -9, -74, -8, 103, 19, -89, 25, 64, -104, 54, -24, -34, 109, -88, -56, 9, 57, 8, 22, -30, -46, 106, 19, -22, -105, -59, 103, 47, 47, -113, -48, 43, -32, 127, -88, 34, 29, -56, 92, -66, -6, 69, -70, -82, -8, 32, 77, 4, 77, -100, 12, 58, -128, 81, 3, -124, 127, 61, -39, 18, -7, -98, 65, -4, -128, 127, 127, -128, -31, 74, -2, -44, -73, 127, 13, -88, 1, -58, -38, 43, 41, -64, 73, 47, -26, 71, -47, -18, -15, -43, -30, 127, 40, -128, -55, 83, -22, 88, 102, -64, 3, -46, -108, 127, 37, -85, 37, 7, 40, -10, -103, -103, 121, 113, -60, -59, 0, 87, 63, -22, -114, -113, 117, 85, -120, 21, 127, -115, -47, 77, 48, -55, -128, -10, 40, 45, 49, 72, -104, -56, 66, -51, 28, -41, 72, 127, -113, -85, 85, -4, -128, 127, 27, -23, 20, -52, 30, -41, 65, -27, -128, 126, 75, -128, 75, 110, -73, -32, -1, 18, 55, 22, 3, -115, 20, 103, -128, -42, -13, 91, 96, -128, 31, 126, 39, -128, -68, 72, 6, -41, 15, 45, 78, -104, -58, 127, 8, -100, -74, 13, 110, -24, -128, 124, 13, 65, -7, -93, 11, -14, -3, 77, 11, 17, 51, -128, 104, -64, -54, 103, -99, -42, 127, -26, -128, 95, 83, 51, -15, -128, -79, 100, -19, -35, -8, 42, 24, -48, 127, -11, -32, -28, -83, 24, -43, 125, 76, -128, 108, 12, -64, 2, -24, 89, -60, 55, -15, -117, 113, 126, -122, 31, 30, -96, -9, -9, 127, -32, -22, 70, -1, -61, 8, 103, -85, 1, 30, -7, 48, -97, 53, -25, -89, 26, 30, 37, 39, 8, -53, -5, -53, 59, -22, -11, -39, -64, 127, 44, -66, -19, -28, -65, 110, -26, -128, 34, 127, 73, -128, 31, 18, -128, 127, 75, -126, 42, -37, -42, 19, 71, 96, -39, -27, -72, -45, 86, 46, -75, -9, -12, 62, 106, -81, -19, 82, -6, -128, 70, 68, -128, 63, 55, -78, -2, 127, -24, 34, -93, -23, 42, -14, 66, 9, -49, 1, -42, 42, 41, -112, 26, 30, -18, -54, -6, -31, 0, 127, -34, -121, 32, 3, 88, 43, -43, -72, 1, 127, 102, -97, -54, -4, -72, 19, -22, 39, 127, -71, -71, 24, 11, 100, 9, 25, -115, -128, -1, 42, 127, -75, -80, 127, -44, -128, 37, 107, -81, 31, 76, -128, -20, -9, 28, 56, -30, 0, 127, -64, -25, 45, -39, 17, -40, 19, 9, 4, 28, -34, 83, -19, -70, 36, -65, 85, 26, -30, -4, -9, -5, 39, 48, -70, 27, 71, -24, 24, -91, -42, -32, 40, 127, -78, -95, -77, 127, 56, -74, -29, 65, 0, -42, -6, 0, 113, -123, -115, 88, 31, 20, 76, -86, -81, 45, -55, -2, 30, -57, 69, 127, -97, -43, 97, 21, 1, 12, 1, -92, -20, -26, -14, -47, 92, 124, -51, 9, 41, -128, -86, 79, 78, -53, 3, -5, -39, 127, -57, 23, -82, -128, 127, -25, 5, 62, -128, 51, 41, 49, -85, 31, 21, -128, 127, 104, -128, -34, 127, -128, 26, 28, -71, 98, -18, -74, 95, -25, -125, 87, -34, -45, 103, 83, -40, -49, -40, 42, -46, 10, 87, -126, 40, 74, -37, 10, -5, 25, -29, -63, 64, 127, -41, -128, 53, 127, -54, -42, -73, 17, 127, -128, 6, 93, -23, -44, 48, -66, -32, 127, -66, -103, -86, -19, 127, 22, -10, -68, 54, 127, -128, -34, 92, 7, -13, -51, -1, -62, 64, 70, -47, 58, -42, -12, -35, -22, -51, -18, 106, -90, -12, 49, -35, 45, 27, -102, 113, 5, -128, 127, 108, -86, -68, 55, -37, -76, -22, 123, 5, 36, 35, -128, 127, -42, -4, 62, -92, 127, 37, -128, 80, 14, -126, 43, 28, 86, -65, -48, 95, -11, -78, 22, 94, 36, -128, 66, 127, -128, 31, -3, -105, 30, 4, -9, 0, -1, 20, 94, 81, 52, -60, 4, -121, 46, 0, -80, 127, -63, -93, 0, 124, -29, 21, 25, 7, 87, -107, 2, -53, -107, 127, -12, -76, -25, -17, 106, -75, 38, 0, 51, 79, -54, 48, -34, -12, 49, -82, -69, -3, -17, 80, 76, -15, -60, -46, 36, -8, 46, -4, -56, -24, -65, 127, 39, -93, -79, 127, 9, -52, -5, -86, 35, 97, 108, -4, -73, 12, -81, 14, 127, -106, -62, 83, -81, -116, 8, 117, 19, 53, -79, -30, 127, -128, -54, 63, -57, 48, -18, 0, -8, -55, 98, 14, -115, 62, 11, 6, 31, -63, 57, -37, 63, -14, -128, -6, 24, 24, 66, 80, -123, 27, 81, -128, 110, -21, -66, 51, -4, 103, 3, 18, -115, -43, 35, -35, -24, 57, -34, 13, -12, 24, 7, -128, 19, 32, 10, 4, 55, 72, 74, -40, -56, -30, 52, 4, -41, -20, 57, -14, -106, 109, -32, -21, 22, 12, -63, 3, 64, -92, 11, 57, -69, -10, 114, -95, 19, 116, -63, -87, 38, 51, -126, -7, -7, 89, 127, -55, -90, 55, -69, 0, 122, -95, 9, -39, -75, 127, -79, -1, 43, -60, 51, -23, -36, -56, 81, 125, 53, -128, -108, 98, 70, -83, 45, 94, -128, 43, 40, -51, 55, -22, -20, -10, -69, -42, 108, 42, -128, 76, 31, -85, 13, 49, 78, -70, 24, -2, -90, 85, 9, -14, -8, -103, 127, -10, -2, 8, -128, 47, 116, 49, 19, -62, -106, -43, 53, 127, -45, -45, 31, -7, 48, 36, -115, -22, 9, -122, 127, 64, -42, -5, -128, 127, 31, -4, -25, -116, 10, -19, 81, 83, 62, -61, -124, -37, 52, 79, 70, 38, -128, -46, 70, -73, -38, 117, 53, -73, 27, 27, -128, -8, 127, -105, -57, 28, 87, 56, -89, -97, 82, -18, -7, 127, -112, 55, 58, -27, -26, -18, 11, 36, -72, -95, -30, 86, -21, 31, 5, 11, 54, -128, 37, 8, -49, 122, 31, -122, 31, -55, -22, 71, -63, -32, 127, 44, -128, 95, 19, -12, 71, -128, 32, 127, -98, 0, 46, -76, 22, 55, -32, -111, -42, -26, 60, 56, 54, 86, -31, -113, 74, -65, -37, 3, -93, 127, 13, -44, -3, 76, -25, -128, 127, -2, -128, 76, 127, 48, -128, 30, 110, -71, 70, 22, -65, -31, -70, 31, 21, 55, 102, -99, -128, 71, 57, -56, -18, 81, 78, -32, 4, -128, 41, 124, -128, 81, 0, -128, 127, -43, 58, 12, -70, 127, -128, -88, 92, -57, 90, 108, -128, 46, 9, -115, 77, 40, 10, 48, -36, -60, 59, -68, 3, 60, 23, 54, -57, -123, -61, 43, 34, -46, 66, -38, 76, 99, -128, -26, 81, -10, -128, 127, -13, -123, 41, 31, 99, 42, -77, -82, -10, 127, -4, -12, 42, -128, 86, -46, -90, 127, -46, -20, -69, 22, 127, -128, -18, 27, -22, 21, -14, 59, -53, -18, 120, -59, 48, 19, 27, -39, -60, 47, -86, -15, 3, 115, 40, -128, 79, 127, 22, -125, -40, -5, -96, 90, -35, 34, 77, -59, 49, 55, -10, 23, -122, -74, 127, 68, -57, -7, 69, -90, -128, -6, 51, 9, 69, 85, -103, -12, 69, -77, 57, -11, -110, 127, 28, -109, -13, 109, 47, -128, 22, 43, 15, 46, -37, 18, -34, -55, 15, 6, 15, 18, -1, -128, 72, 57, -40, 0, -128, 39, 80, 66, -14, 2, 52, -128, -66, 43, -53, 127, 24, -36, 27, -109, 49, -6, -80, -11, 100, 81, -11, -40, -45, -11, 27, -18, 56, -13, -48, 99, 14, -126, 15, 39, -117, 40, 66, -35, 40, 44, -54, -79, 12, 127, -39, 22, 120, -93, -128, 75, -8, 31, -9, -43, 18, -12, 126, 25, 3, -85, -20, 20, -13, -44, 31, 52, -8, -96, 60, 21, -45, 0, -51, -34, 100, 92, -21, 61, -128, -128, 105, 2, 53, 55, -46, 98, -121, -66, 126, 75, -128, -73, 107, -19, 65, -56, -109, 59, 42, -92, 92, -9, -86, 34, -37, 11, 94, 127, 24, -24, -128, -53, 127, 75, -128, -19, 127, -123, -92, 123, -40, -54, 8, 38, 114, 25, 12, -128, -60, 57, -53, -8, 20, 47, -19, -18, 48, 103, -52, -71, 83, -55, 59, 61, -128, 99, -5, 21, -28, -92, 127, -100, 41, 102, -30, -5, -17, -14, 32, -117, 14, 127, -128, -119, 26, 39, 3, 74, -49, -42, 127, -14, -65, 87, -128, 4, 127, -128, 23, 73, -2, -72, 15, 66, -128, 34, 24, 24, -21, 29, 90, -12, 1, -40, 47, 18, -128, -93, 98, -55, 52, 51, -25, 17, -87, 71, -22, 23, 119, -8, -60, -34, -41, -37, 5, -37, 127, -13, 19, -37, -128, 127, -48, -126, 121, -27, 54, 107, -124, -39, 58, 107, 1, -122, -58, 110, 91, -88, -24, 59, -57, -78, -1, 62, 34, -40, 60, -19, -9, 69, -55, -108, -1, 93, -49, -115, 113, -6, -2, -15, -42, 88, -93, -31, 121, 31, -117, 70, -53, 54, 85, -100, -29, 90, -44, 6, 81, -128, 30, 73, -91, -51, 127, 52, 40, -119, -19, 127, -119, -23, 90, 63, -128, 45, 21, -46, 71, -89, 15, 23, -36, 71, 106, -77, 3, -88, -26, 48, -59, -35, 96, 32, -96, 65, -60, -49, 102, 107, -128, 31, 73, -43, 90, -97, 32, -77, -95, 73, -4, 71, 52, -9, -19, 8, -47, -13, -69, -102, 127, 17, -128, 102, 51, -13, -70, 34, -36, -128, 127, 13, -126, 43, -18, 117, 127, -128, -100, 39, 49, 40, 105, -55, -120, 127, -81, 34, 70, -128, -31, 45, 69, 7, -48, -20, -3, 76, -25, -66, 112, 78, -58, 17, -77, -32, 127, 20, -27, -18, 54, 49, -128, 12, -2, -63, 97, -74, -31, 127, -35, -70, -10, 39, 116, -71, -128, -31, 11, -5, 49, 83, 66, 22, -98, 29, 15, -128, 60, 127, 11, -81, 46, -88, -62, 11, 47, -9, -56, 52, -96, 109, 123, -113, -5, 56, 11, 1, -14, 18, 22, -128, -42, 96, 47, 42, -71, -81, -71, -4, 32, 98, 97, -116, -128, 40, 54, 66, -12, 34, -81, -64, 127, 43, -128, -55, 106, 57, -60, -93, 125, -74, -21, 38, 28, 57, -103, -31, 127, -29, -42, 8, -76, 60, 46, -24, -94, -40, 43, 88, -49, -26, 15, 89, 9, -124, 27, 122, -74, -26, 26, 18, 82, -5, -102, -32, 58, -49, 123, -43, -30, 70, -32, -76, -53, 23, 57, 3, -56, 98, 80, -75, -128, 127, 3, -113, 10, 37, 7, -94, 127, -13, -38, 85, -18, 76, -128, -102, 31, 127, 0, 0, 4, 11, -88, -41, 35, -62, 127, -31, -117, 43, 83, -63, -43, 97, 3, -39, -56, 12, 88, -96, 46, 38, -9, 63, -106, 41, 105, -80, 14, -44, -41, 26, -60, 31, 127, -70, 5, 80, -61, -86, -59, 32, 8, 45, 87, 43, -128, -115, 62, 91, -62, 69, 124, -44, -29, -128, 41, 38, -10, 12, 3, -55, 7, 127, -32, -13, -91, 15, 34, 8, 76, -30, -116, -59, 20, 127, 127, -128, 47, -4, -46, 12, -120, 87, 126, -3, -51, 9, -111, -56, 127, 37, -119, 30, 15, -108, -14, 87, 54, 11, -61, -14, -11, -21, 71, 2, -47, 15, 58, -47, 21, 8, -65, 86, 86, -97, -64, 40, 71, -30, -22, 94, -128, -96, 93, 36, -58, 76, -72, 39, 78, -128, 22, 30, 71, -107, -107, 29, 66, 96, -23, -64, -81, 127, -27, 13, 38, -90, 87, -78, -72, 32, 127, -68, -65, 79, -28, 97, -82, -53, 127, -1, -128, -32, 39, 80, 9, -109, 105, 105, -128, -64, 42, -61, 34, 25, -48, 42, 124, -6, -38, 40, 58, -60, 12, 20, -128, 31, 82, -55, -26, 30, -46, -18, 127, -13, -91, -35, 107, 7, -128, 127, 85, -107, -122, 126, 98, -128, 12, 32, 42, -35, -105, 108, 96, -94, -89, 127, 79, -12, -86, -93, 23, 25, 38, 126, 5, -24, -72, -34, -13, -23, 57, 43, 53, -74, 14, -37, -20, -19, 6, 20, -86, 89, 82, 7, -14, 21, -26, -81, 14, 45, -24, -1, 64, 40, -38, -75, 22, 48, 36, 1, -128, -49, 52, 77, 25, 27, 37, -4, 35, -113, -128, 127, 116, -90, -5, -43, -62, 125, 20, -49, -25, 34, -23, -128, 86, 91, -34, -86, -1, 8, 74, 13, -81, 124, 80, -26, -10, -30, 7, 29, -128, 40, 127, -52, -18, -58, -90, 114, 21, -59, 58, 3, -25, -1, 81, -128, -52, 52, -68, 95, 21, 3, 98, -31, -34, 29, -19, -43, 5, -2, -45, 25, 31, -98, 21, -17, 0, 115, -99, -120, 62, 112, 68, -128, -30, 127, -104, -123, 127, 11, -37, 39, -128, 105, -28, 30, 92, -43, 19, -90, -1, -24, -53, 3, 38, 114, -19, -115, 45, 73, -55, -88, 44, 13, -51, -25, 127, 28, -128, 123, 42, 27, -77, -42, 124, -104, 19, 27, -98, 6, 100, 44, -19, -128, 93, 7, -28, 66, -106, 54, -80, 38, 111, -76, 51, 49, -75, 30, -109, 3, 105, -55, 25, 29, -66, -38, -26, -78, 127, 19, -78, 94, -81, -96, 127, -31, -77, 111, 0, 41, -72, -32, 71, 40, -77, -61, 97, 44, -74, -1, 42, 31, -24, -115, 71, 65, -3, 0, 18, -12, -128, -14, 48, -53, 76, -41, -37, -11, 76, -39, -2, 127, -82, -86, 40, 71, -128, -41, 122, -40, -48, -14, 1, 80, 52, -123, 4, 51, 69, 17, -128, -51, 127, 54, -106, 44, 18, 36, 25, -100, 36, 51, -100, 0, -32, -48, 41, -28, 59, 119, -37, -128, -80, 127, 78, -73, 69, -78, -128, 127, 97, -128, 92, 61, -69, 12, -80, -5, 56, -87, 93, 48, -28, 24, -128, -51, 127, 51, -86, 35, 23, -116, 45, 88, 38, -34, -128, 114, 41, -114, 65, -44, -42, 110, 22, -76, -97, 127, 58, -47, -102, 6, 3, 65, -11, -123, 11, 90, 111, -85, -28, -53, 32, -30, 45, 70, -102, 127, -55, -10, 20, -20, 127, -34, -66, 4, -108, 29, 103, -38, -23, 7, -37, -13, 71, -81, 45, 72, -128, 11, -4, -19, 109, -14, -13, -41, 55, 106, -128, 48, 85, -116, 60, 23, -106, 0, -3, -13, -12, 110, -59, -30, 111, -95, -8, -43, 61, -7, 1, 100, -42, 27, -80, -79, 17, 63, 24, 71, -26, -70, 109, 59, -128, -13, 90, -64, -54, 58, 104, -74, -26, 85, -78, -99, 0, 71, 5, 18, 95, -128, -26, 58, 29, 38, -27, -110, -43, 2, 119, 75, -73, 74, -52, 1, 49, -128, -19, -1, -76, 57, 81, 83, -91, 52, -26, -86, 116, -18, -30, -12, 64, -107, 55, 89, -61, 25, -53, 77, 18, -92, 2, -14, -15, -42, -2, 6, -25, 127, -39, -65, -14, 86, 7, -100, 127, -55, 40, 13, -24, -2, 6, 34, -103, 55, 126, -128, -107, 121, -87, 74, 127, -90, -94, -25, 63, 44, -24, -117, -9, 127, -41, -26, 25, -31, 93, -76, -38, 123, -55, -69, 126, -55, -27, 17, 6, 91, -113, -63, -12, 32, 4, -56, 127, 51, -87, 47, -48, -106, 89, 86, 19, -110, -87, 46, 52, -38, -18, 11, 53, 109, -62, -17, 94, -63, -128, 127, -7, -100, 45, -47, 121, 1, -68, 68, 54, 61, -85, -128, 0, -26, 109, 127, -128, -128, 27, 105, -24, -29, 110, 55, -83, -103, 82, -20, -6, 82, -102, -4, 127, -104, -17, 87, -61, -57, -32, 41, -27, 44, 51, -73, 49, 1, -92, 102, 10, -65, 13, -7, 82, 115, -111, -128, 19, 127, -22, 8, 17, -83, 36, -42, 51, -24, 15, 127, -128, 18, 15, -114, 57, 36, 0, 62, 31, -60, -31, 48, 52, -27, -117, -9, 93, -70, -10, 110, -128, 10, 109, -113, -74, 114, 31, -72, 122, -114, -45, 35, -127, 127, 65, -72, -25, 106, 17, -128, 52, 127, -128, -74, 127, -59, -86, 32, 65, 87, -91, -21, 87, 20, -104, -128, 127, 81, -54, 34, 15, -107, 34, 111, -128, -41, 40, -3, 24, 26, 40, -119, 25, 97, -8, -46, 47, 86, -24, -43, 21, -75, -63, 120, -81, -8, 127, -128, -68, 79, 97, -96, -21, 127, -128, -128, 90, 29, -1, 75, 55, 27, -14, -81, -20, -20, 63, 21, -120, 82, -19, -87, -24, 117, -11, -100, 127, -105, 5, 28, -15, 97, -64, -2, 39, -37, -4, 86, 23, -128, 10, 119, -128, 6, 9, 4, 127, 66, -128, -128, 127, 5, -76, 127, -73, -43, 23, 35, 71, -128, -77, 61, 86, 3, 56, -70, 5, 79, -128, 40, 64, 30, -73, -24, 26, -60, 10, -25, 17, 31, 27, -55, 48, 127, 26, 6, -72, -98, 87, -31, -106, 127, 22, -128, 13, 81, -53, -19, 127, -36, 9, 39, -128, -18, -15, 34, 69, -45, 6, 80, -19, 23, 52, -128, 9, 119, -124, -52, -7, 126, 61, -116, 90, 86, -77, -92, -10, 61, 66, -74, -115, 83, 124, -122, 24, 102, -55, -102, 60, 127, -31, -117, 10, 21, -58, 17, -77, 17, 107, -87, -47, 127, 12, -128, 78, 127, -68, -128, 48, 5, -44, 78, 87, -117, 1, 102, -10, -60, 1, 81, -115, 12, -32, -95, 7, 71, 72, -110, 87, 127, -128, -121, 127, 36, -95, 43, -14, 31, 59, -9, 70, -128, -77, 127, -75, -77, 43, 110, 41, -128, 12, 122, 7, -21, -128, 59, 43, -128, 127, -66, -128, 127, -45, 10, 38, -97, 42, 25, -32, -86, 64, 0, -34, -53, 127, 75, -128, 21, 2, 93, 54, -128, 73, 68, -47, 87, -69, -128, -1, 71, -58, 41, 35, -55, 46, 37, 69, -110, -78, 42, -37, 127, 2, -78, 115, -64, 41, -36, -40, 74, -127, 20, 86, -60, -94, 86, -5, 0, 86, -47, 65, 55, -128, -44, 6, 35, 127, 31, -42, -94, -113, 127, -6, -99, 73, 71, 57, -85, -106, 23, 127, -51, -128, 49, 85, -95, 96, 73, -68, 19, -125, 42, 43, -128, 127, 6, -62, 126, -106, -99, 127, -31, -128, 127, 47, -112, 107, -77, -1, 127, -59, -10, -97, 27, -5, -44, 127, -110, -113, 92, 63, -49, -95, 114, 37, -128, -58, 127, 122, -128, -83, 125, -10, -75, 83, 42, 32, -47, 9, 59, -94, -2, 12, 8, -18, 12, 0, -87, 99, 68, -128, 21, 19, -89, 95, 28, -51, 30, 6, 77, 37, -82, 9, 28, 58, -107, -70, 94, 37, -66, -28, -11, -62, -43, 127, 63, -32, -36, 17, 97, -128, 64, 70, -128, -25, 127, 48, -85, -30, 96, 20, -128, 61, -5, 47, 76, -106, 9, -12, -58, 100, 107, -111, 30, 90, -114, -51, 59, 42, -36, -64, 86, -19, 15, -82, -39, 127, -30, -92, -70, 75, 81, -63, -96, 125, -25, -13, 15, -46, 127, -53, -100, 74, 66, -79, -13, -40, 64, 0, 11, 22, -57, 93, 9, -47, 10, 1, -87, -9, 62, 25, -126, -34, 127, -42, -102, -51, 127, 55, -100, 98, 42, -128, -9, 115, -57, -68, 85, 0, -60, 90, 25, -86, -4, 78, -128, 18, 48, -23, 1, -68, 12, 29, 85, -62, -2, 127, -124, -18, 29, 4, 74, -128, 69, 14, -23, 4, -45, 55, 6, -75, -36, 43, -3, 108, 78, -104, -31, -56, 68, 111, -128, -72, -42, 127, 5, -46, 117, -78, -38, -39, -24, 0, 11, 3, -11, 127, -39, -22, 36, -25, 80, -10, -128, -68, 104, 92, 10, -125, -106, 86, 127, -87, -30, 127, -128, 19, 79, -14, -22, -128, 127, 93, -128, -35, 99, 26, -96, 109, -6, -57, 114, -110, -56, 127, -32, 40, 65, -128, -78, 117, 69, 22, 63, -125, 9, -31, -98, 62, 114, 24, -124, 105, -70, -71, 25, 1, 127, -76, -81, 127, 83, -128, -117, 31, 119, 34, -119, 5, 62, -55, 117, -26, -128, 127, 7, -18, 109, -59, -119, 77, -32, -45, 127, -92, -120, 127, 92, 7, -102, -128, 127, 127, -128, 26, -22, 5, 51, -128, 9, 78, 32, -108, 57, 72, -122, -75, 59, 127, 9, -60, 28, 15, -75, -54, 120, -15, -116, 71, -2, -64, 120, -52, -69, 6, -60, 107, -26, -36, 127, -27, -111, 0, 97, -97, 44, 127, -128, -48, 119, 55, -121, -30, 82, -42, 103, -30, -13, 12, -128, -6, 108, 122, -65, -115, -55, 70, 127, -88, -120, 105, 75, -52, -87, -5, 41, 127, -79, -94, 81, 45, -44, -31, 11, 1, 127, -86, -128, 127, 80, -128, -64, 47, -2, 27, 77, -64, -54, 27, 43, -28, 91, 116, -91, 36, -89, -5, 127, -128, -63, 28, 78, 31, -9, -68, -111, 127, 0, -93, 51, 91, -40, -57, 127, -54, 1, 18, -112, 127, -2, -36, -60, -56, 81, 43, -63, -1, 74, -117, 30, 127, -95, -44, 0, 91, 28, -113, 41, 29, 9, -103, -57, 127, 18, -116, -32, 25, 55, 41, -77, 102, -4, -128, 42, 45, 94, -30, -110, -15, 42, 106, -98, -3, 51, -93, 85, 43, 14, -73, -66, 31, -22, 62, -36, 5, 126, -80, -122, -1, 127, -15, -128, 127, 28, -96, 46, -21, -122, 95, 107, -80, 5, 52, -95, 62, -46, -3, 100, -24, -83, 39, 0, -100, 97, -34, -58, 1, 85, -38, -1, 46, -53, 89, -31, 25, -18, 21, -3, -128, 116, 69, 5, -78, -24, -45, -52, 127, -93, 58, 97, -128, 96, 60, -44, -40, 37, 75, -45, -73, 81, -58, -24, 60, -128, -7, 49, 25, -26, 19, 74, 78, -70, -65, 6, 63, 34, -47, -3, -14, 5, 57, 35, -98, -22, -6, 52, 7, -110, 11, 127, -72, -35, 103, -43, -3, 45, 37, -128, -125, 59, 127, -91, 0, 57, -78, 57, 94, -94, -128, 86, 103, -79, -57, 13, 52, 120, -128, -80, 10, 77, 4, -51, 35, 111, -62, -128, 127, 127, -109, -128, 46, 21, -48, 4, 65

	
	);
 
    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project
 
    constant SCENARIO_ADDRESS : integer := 0;    -- This value may arbitrarily change
 
    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
 
                o_done : out std_logic;
 
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;
 
begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
 
                o_done => tb_done,
 
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );
 
    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;
 
    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
 
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
 
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;
 
        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
 
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;
 
        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';
 
        -- Wait some time for the component to reset...
        wait for 50 ns;
 
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
 
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock
 
 
        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
 
        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
 
        wait until falling_edge(tb_clk);
 
        memory_control <= '1';  -- Memory controlled by the component
 
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
 
        tb_start <= '1';
 
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        wait for 5 ns;
 
        tb_start <= '0';
 
        wait;
 
    end process;
 
    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin
 
        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';
 
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
 
        wait until rising_edge(tb_start);
 
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;
 
        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(signed(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;
 
        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);
 
        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;
 
end architecture;

