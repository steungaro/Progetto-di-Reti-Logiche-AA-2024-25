-- TB EXAMPLE PFRL 2024-2025 -- RUAN HUIJUN
 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
 
entity tb2425 is
end tb2425;
 
architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
 
    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");
 
    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 32759;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      126,                                                        -- S
                                                      0, -1, 8, 3, -8, 1, 0, 1, -9, 45, 0, -45, 9, -1           -- C1-C14
                                                      );
    signal scenario_input : scenario_type := (61, 18, 51, 28, -47, -128, 36, -119, -65, -6, -82, 60, 63, 127, -5, -118, -11, -119, 65, -30, 89, -88, 87, 127, -89, 67, 45, 20, -48, 32, 118, -115, -77, 42, 41, 4, 42, -50, 13, 105, 72, 59, 38, 7, 59, -95, 17, -80, -86, -46, 19, -125, -5, -22, -126, 34, -83, 47, -74, -3, -48, -84, 10, 3, 86, -76, -121, 0, 2, 20, -22, -54, -49, -112, 81, -118, -79, -30, -69, -37, 53, 78, -33, -80, -72, -31, 82, -27, -111, -120, 99, -31, -76, -19, 100, -117, 33, 107, 11, -93, -1, 117, -19, 78, -123, -66, 89, -74, 33, -108, 18, -42, 98, 113, 6, -102, -46, -40, -1, -29, -32, -30, 68, 20, 80, 40, 31, -15, 19, -85, 21, -110, -96, -126, 97, -90, -63, 58, -36, 98, 78, 110, -72, 48, 95, 62, 74, -78, -106, -55, 21, -10, 44, -38, -118, -4, -126, 42, 109, 22, 85, 2, 40, 117, 5, 9, -101, 70, -61, -8, 40, -111, -26, 96, 65, -58, 30, 11, -8, 52, 85, -115, -86, 1, -25, -76, 125, -22, 94, 106, -128, 51, -19, 40, 41, 114, -78, 68, 56, -11, -68, -32, 7, 35, -64, -56, 105, 94, 84, -31, 18, 41, -18, 60, -86, 86, 112, -89, -64, 79, -111, -64, 2, -2, 104, -85, -16, -102, 112, -88, 16, -84, 8, -105, 79, 72, -33, 56, 38, -77, -103, -72, 92, 8, 116, -122, -34, 101, -83, 30, 52, -65, 94, -74, 61, 70, -30, -82, 97, -46, -42, -15, -2, 95, 8, -50, 39, 103, -122, -50, -101, -96, 6, 119, 40, -5, 126, -122, -32, -85, 36, -108, -22, 2, -54, -88, -56, 44, -42, -87, 126, 44, 26, -3, 11, -94, 75, -77, -118, 81, 1, -91, 113, -121, -100, 25, 2, -102, 31, 98, -58, -61, 118, 48, 69, -63, 88, -114, 109, -82, -73, 108, 91, 82, -23, -26, 116, -76, 25, 126, -123, -102, -93, 119, -94, -64, 16, 36, -38, -80, 7, 32, -13, -3, -47, -71, 62, -87, -57, 44, -40, -2, 24, -77, -48, -127, 25, -59, -75, -77, -61, -70, -51, -25, -79, -17, 39, 66, -108, -127, 114, 27, 34, -27, -104, 115, 30, 87, -100, 101, 3, -12, -28, -101, 39, 52, -100, -63, 121, -47, -12, -67, 11, 65, 36, 61, -79, -53, -1, -59, -52, -15, 96, 110, 86, 120, 97, -11, 79, 126, -38, -46, -14, 62, -19, -102, -13, 9, -37, -20, 90, 79, 41, -26, 16, -51, -93, 65, 24, 34, -122, 101, -109, 102, 83, 105, 95, 53, -34, 46, 51, 57, -127, -91, -9, -18, -65, 106, 120, 26, -41, 82, -23, -128, -72, 122, -50, -37, 59, 102, 125, 66, 75, -112, 40, 31, 122, 7, -44, -40, -74, -121, -111, -73, -84, 9, 37, -20, -13, 29, -122, 74, -16, -16, 75, 40, -22, -103, -124, -91, 127, -127, 103, 75, -110, 16, -22, -116, -105, 62, -28, -51, 69, -10, 4, 113, 127, -86, -35, -14, 71, -28, -67, -73, 84, -120, 96, -66, -95, 100, -29, -96, 101, -53, 107, 119, 91, -43, -125, 114, -109, -24, -64, 88, 94, 68, 74, 93, 110, -89, -49, 54, 11, 12, 109, -33, 20, 77, 29, 53, 49, -127, 86, 23, -52, 65, 14, -89, -105, 18, -103, -86, 122, -39, -125, 88, -98, 77, 53, -116, 116, -124, 66, 0, 17, 48, 95, -91, -3, -3, 91, -81, -2, 49, 70, 74, -14, -44, 113, 9, 102, -118, 52, 96, -28, 55, 56, 2, 4, -19, 14, -8, -14, -47, 120, -125, -127, 88, -88, -2, -43, -125, 45, 83, 52, -13, 29, -89, 72, 14, 48, 46, 24, -28, 15, 124, -101, -57, -2, 31, 53, -115, -104, -89, -34, -112, -86, -33, 104, -46, 93, -67, -42, 11, -112, -118, 126, 45, -79, 70, -69, 98, -11, 84, -58, -124, 80, -30, -53, -49, -127, -128, -36, -103, -89, 58, -86, -47, -103, -110, 36, 118, -48, 122, 1, -32, -124, 0, -114, -74, -58, -55, -104, 59, -99, -34, 63, 110, 64, -117, -67, 66, -117, 25, 91, -77, -45, -123, 4, -20, -104, -88, -30, -24, -94, 100, 72, -89, -28, 86, -35, 42, -96, -11, -26, -67, 83, -91, -85, 20, -80, -24, -42, -68, -127, -79, -17, -44, -73, 115, 64, -49, -100, -93, 55, -66, -121, -1, -27, -21, -42, 66, -107, -10, -73, -5, 51, -117, 33, 95, 31, 81, -57, 117, -115, -55, -90, -4, 29, -35, -16, -34, 44, 12, 1, -29, 74, 8, 99, -80, 115, -71, 114, -120, 47, -86, 4, -30, -75, -91, -63, 84, 118, 9, 73, -124, 82, 111, 0, -17, -51, 112, 77, 121, -4, -50, -35, -57, 86, -64, -9, 73, -7, -23, 82, -88, 19, -42, 10, 72, -5, 76, 28, -15, -43, -27, -11, -89, -43, 118, 22, 34, 102, -28, 27, -29, 50, 120, 42, 9, -72, -95, -46, 49, 10, -92, 89, -98, -6, -28, 102, 117, -80, 3, -25, 5, 104, 92, 44, -67, 82, -62, 95, 57, 38, -5, -100, -39, -13, 70, 98, 44, 103, -76, -35, -15, -39, -73, 15, 83, 27, -10, 73, 75, 121, -80, -48, 97, -116, 124, -97, 95, -66, 126, 24, 101, -7, 52, -66, 109, -6, -96, 25, -31, -44, 118, 82, 45, -83, -30, 1, 72, 88, -54, 19, 81, -6, 99, 50, 6, 95, 81, -27, -98, 80, 125, -125, -55, 49, -63, -74, -85, -31, 79, 12, 53, 70, -33, -29, 115, 65, 100, 60, 25, -82, -49, -22, 40, -77, -100, -82, -110, 110, 20, -80, 62, 17, -77, -121, -61, -12, -66, -18, 85, -115, 123, 11, 83, -38, 110, 71, -101, 82, 3, 52, -128, 82, -98, 40, -123, -70, 86, -104, -88, -22, -56, 102, 124, -4, 110, -65, 112, -84, 45, 70, -71, 40, -47, -115, -126, -65, 84, -99, -111, -41, 81, -111, -87, 111, 57, -81, -86, 15, -57, -46, 122, 15, -71, 118, -117, -89, -75, 124, -45, 98, 66, 12, 11, -109, 25, 13, -46, -19, 43, -29, 68, -4, -12, 110, -20, -83, -99, 22, 60, -28, 104, 54, 115, -95, 44, 127, -56, 97, 123, 27, 68, 61, -88, -49, 80, 65, 92, -94, -81, 7, 5, 115, -124, 121, 97, -16, -90, 126, -122, 98, -30, 110, 25, -42, -112, -59, -43, -40, -89, -48, 116, 107, -115, -100, -70, 93, 93, -106, 127, -116, 30, 4, -128, 34, -3, 97, -110, 35, 96, -104, 5, -62, -122, -98, 24, -106, -28, 109, -17, 11, -67, -29, -10, -54, -1, 48, -89, -36, 70, -90, -23, -28, 42, -23, -122, -89, -54, -104, 74, -86, -80, -48, -19, -73, -18, -123, -51, 82, 115, 60, -35, -80, -97, 83, -5, 30, 3, 34, 123, -54, 73, -28, 46, -13, 77, 53, 27, -105, 77, -27, -62, 126, 53, 47, -75, -92, 52, 2, 118, 39, -65, -44, 88, -34, -89, -45, 125, 43, 117, 120, 117, 62, -36, 35, -78, -87, -40, 77, -64, -90, -78, 2, -92, 104, -79, -39, -116, 102, 91, -126, 13, -102, -42, -27, -7, -2, 56, -10, -87, 46, -18, -98, -20, 74, 65, 30, 115, -102, -21, -77, -64, 30, 54, -28, 6, 103, 61, 18, 77, 24, 20, -37, 51, 107, 64, -84, -23, -7, 34, 18, -89, -112, 48, 19, 90, -15, -78, 77, 11, 29, -128, 75, -69, 54, -81, 65, 30, 108, -45, -21, 5, 104, 70, -72, 83, 7, -28, -68, -128, -122, 78, -89, -106, -2, 58, 112, 111, 108, 61, -5, 10, 61, -58, 69, -12, -10, 7, -110, -30, 90, -3, 103, 66, -60, -97, 21, 75, 3, 81, 75, 9, 31, 114, 31, -99, 44, 15, -115, 25, -52, 8, -93, -118, 78, 104, -2, -60, -17, 16, 39, -54, -115, 14, -116, -47, 46, 34, -100, -79, -13, 103, 59, -109, 89, -38, -80, 6, 106, -67, -97, -74, 69, -62, -64, 20, -86, 62, 88, 26, -50, -1, 100, -36, -114, 112, 45, 60, 18, 74, 109, -122, 49, 40, -103, 11, -125, -55, -111, 109, 7, -80, -93, -52, -14, -28, 96, 28, -94, 57, -74, -15, -72, -102, 77, -58, -117, -6, -126, 29, -60, 112, 35, 118, 24, 60, 1, 27, -122, 18, 8, 13, 66, 44, 89, -76, -112, 58, 80, -78, -13, -121, 35, 43, -95, -16, 114, -84, 107, 116, 74, -81, 100, -19, -91, -3, -86, 38, -104, -80, -72, 33, 61, 122, -51, 22, -82, -35, -48, 127, 15, 67, -122, -77, -17, -89, 35, -31, -44, 14, -43, -98, 62, -70, 11, 99, 55, 53, 10, 79, 101, 66, -16, 34, 61, 61, -71, 107, -102, 9, 106, 42, -51, 112, 93, 60, -104, 0, -99, -20, -113, -14, 10, 77, 44, -107, 48, -29, 75, -70, -77, 48, 125, 35, -45, 58, -31, 12, 37, -5, -107, 16, -91, -30, 0, -126, -98, 24, 3, -69, -124, 18, 46, 14, -33, -38, 36, -113, 62, -17, -54, 113, -97, -57, 20, -14, -127, 117, 126, 38, -15, -108, -74, 22, -10, 55, 25, 21, -49, -100, 80, -44, 46, -2, 98, -115, 89, 6, -100, 23, 117, -26, 8, -107, 45, -100, 7, 46, -110, 6, -43, 3, 26, 11, -103, -112, -62, 50, 37, 18, 78, -10, 102, -4, 116, 72, 9, 77, -49, 38, -28, -60, -116, 108, -39, 58, -119, 97, -24, -101, -25, 61, 30, -127, -55, 55, -111, 11, -22, 55, -99, -72, -83, -125, 53, -95, 76, -66, 111, -101, 100, -45, -33, 113, -64, 57, 43, -55, 26, -109, -28, -127, 81, -126, -126, -102, 57, -109, 37, -93, 74, 67, -36, 119, 70, -111, -103, 18, -49, -120, 45, -76, -37, -115, -91, 27, 70, 80, 100, -32, 99, -56, -31, 52, -54, -29, 78, -124, -10, -12, -89, -63, -73, 3, -72, 125, 20, -47, 16, 100, -39, -67, -104, 53, -54, -67, -48, -112, -115, -75, -16, 112, -3, 81, 37, 72, -76, -13, 76, 43, 103, 115, 108, -98, -9, -92, -100, -117, -10, 44, 111, 79, 105, -121, 4, -76, -60, 85, -60, -47, -118, 53, -62, 7, 6, 103, -49, 59, -38, -101, -26, -62, -113, -46, -32, 6, -10, -4, 17, 108, -88, 1, 60, -110, 8, -64, -58, 77, -107, 10, -98, -97, -65, -32, 39, 70, -57, 118, 1, 34, -110, 103, 100, -95, -71, -60, 39, 47, 65, -72, 28, 105, 57, -40, 123, -62, 24, -63, -113, 46, 76, -83, 77, -117, 14, -12, 81, 85, -21, -46, -9, -3, -71, -37, 30, -14, 32, -59, -94, -31, -3, 62, -54, -73, -106, -58, -7, 46, 7, 8, -36, -45, 53, -86, -33, -61, 30, -80, -103, -119, 3, 16, 6, 60, 108, -92, -81, 12, -23, -47, 109, 103, -113, -73, -98, -91, -3, 23, 83, -123, -97, -80, -40, 84, -38, 55, -104, 120, 104, -79, -126, -21, 65, 8, -89, 45, 45, -42, -71, -106, 39, -90, 125, 54, -34, -101, 91, 91, 50, 47, 96, 81, 95, -71, 38, -71, 112, 62, -79, 88, 111, -77, -61, 48, 60, -21, -34, -23, 65, 23, -1, -23, 62, -3, -97, -100, 24, 123, 119, -53, 42, 88, -100, 9, -111, 66, 66, -127, 0, 115, 90, -17, -89, -99, -96, 99, 8, -2, -52, -54, -107, 75, 51, 83, -56, 82, 111, 97, 77, 103, -84, -9, 63, -56, -128, 80, -117, 66, 81, 11, 54, 43, 123, 93, 73, -101, 64, -47, 25, -116, 27, 46, 87, -50, 2, -96, -95, -15, -127, 110, -40, -83, -26, -105, -11, -26, 103, 0, -87, 57, -116, 95, -28, -121, 60, -83, -94, -4, -1, 59, 8, -102, -23, -33, -23, 107, -1, 10, -35, 0, -8, 53, 45, 94, 77, -93, -59, 52, 35, -18, -19, 47, -51, 82, 54, -119, 127, 88, 5, -2, 19, -115, 25, 125, -20, -126, 104, 108, 12, -59, -20, -124, 123, -102, 99, 72, -67, -88, -4, 96, 22, 106, 16, 99, 60, -58, 108, 59, -97, -15, -70, 50, -2, 83, 47, 106, 85, 24, 86, -31, 93, -61, -27, 88, -35, -56, 32, 26, -16, -99, -6, -122, -121, -118, 105, 67, -47, 85, -2, -16, -58, 56, -94, 68, 11, 82, 47, -32, -22, 5, 65, -57, 72, -89, -96, -91, -17, 64, 63, 96, 93, -70, 102, 100, -60, 80, 39, 21, 37, -90, -123, 108, 94, -88, 48, -22, 122, -33, 74, -28, 101, 12, 43, 45, 51, 75, 83, -94, 12, 18, -126, -23, 76, 105, -50, -111, 57, 117, 38, -34, -101, 44, -54, 122, 84, 123, -28, 78, -38, -82, -78, -65, 58, 93, 109, -19, 41, 64, 16, -75, -46, 18, 30, -97, -5, 108, -80, -76, 98, 86, 19, 125, 2, 93, 119, -42, 88, -37, -92, -77, 10, -42, -14, -60, -76, -33, 50, 93, -97, -62, -110, -14, 84, 48, 17, -48, 29, 65, 4, -1, 23, -105, -4, -102, 117, -12, -16, 77, 79, 21, -128, -39, 107, -13, 30, -97, 82, -48, 124, 114, 18, -114, -28, -26, 63, 117, 54, -36, 54, -69, 91, -51, -46, -41, -25, -57, 75, 88, -107, 27, -19, -107, 116, -40, 8, 18, -8, -37, 98, -12, -51, -12, 3, 49, 91, -62, 38, 17, 30, -36, 76, -7, 41, -97, 80, -111, -26, 28, 105, -5, -73, -42, 17, -85, 46, -103, 62, -90, -12, 32, 27, 65, -107, -98, -14, 112, -32, -104, 1, 126, -12, -50, -9, -98, -19, -57, -81, 83, 99, -104, -49, -102, -18, 96, -58, -100, 121, -124, -61, -18, 36, 94, -81, 57, 124, 34, 41, -36, 58, -85, -38, -81, -7, 81, -51, 102, -104, -4, 57, 124, 20, -120, -106, -126, 104, -36, -98, 98, -32, -31, -48, -123, -65, -1, 62, -69, -95, -24, 23, 92, 19, 113, -117, -116, 66, -40, 114, 91, 84, 43, 87, -24, 52, 109, -22, 28, -54, 8, -2, 42, 106, 78, 47, -87, -50, -18, -27, -17, 86, 124, -53, -23, 110, -42, -11, 48, 46, -25, 11, 2, -110, -30, 106, 70, -48, -44, -29, 26, 93, 97, -60, 71, 48, 116, 112, 126, -30, -43, -19, -72, -46, 57, 33, -64, -113, -106, 112, 62, -3, -4, -64, 15, 94, -85, -42, -82, -1, 57, 72, -36, 26, -115, -93, -54, -127, -108, -56, -29, -23, 54, 27, 59, -17, -68, 123, -2, -46, 108, -68, 79, -24, -3, -34, -58, 40, 52, -11, -89, -19, -67, 4, -120, -54, 39, -46, -53, 59, 27, 46, -91, -47, -55, 96, 64, 5, 92, -66, 87, 72, -5, 38, -80, 120, -123, -10, 32, 57, 107, 71, -89, -87, -53, -81, -13, 115, 1, 63, 46, -100, -19, 83, -19, 55, 52, -83, -68, 16, -20, -108, -40, 103, 58, 8, 95, 63, 126, -1, -7, 106, -58, 32, -109, 18, 79, 6, 5, -48, -59, -77, -19, 51, -121, 90, -22, 59, -120, 38, -53, -12, 58, 35, -37, -11, -85, -70, -76, -87, 57, 45, -109, 127, -51, -90, 17, -100, 45, -106, -19, 114, -54, 90, 37, -47, 52, -113, -116, 60, 54, -41, -80, -16, 122, 11, 101, -91, 69, -102, -50, -2, 71, -30, -2, -107, 8, -113, -79, -75, -90, 30, -88, -16, -8, 77, 65, -83, 93, 77, 105, 19, -92, -102, -125, -98, 37, 105, -61, -21, -125, 17, 105, 74, 115, -25, 95, -4, -9, -111, 49, 29, 47, 89, -115, -88, 39, 78, -43, 4, 27, -66, -105, 63, -40, -102, 93, 126, -125, -96, -23, -122, 49, -46, 81, 37, 58, 48, -95, -79, 65, 82, 78, -15, 44, 91, 25, -45, 41, 110, 87, -60, -84, 110, -125, 5, -120, 96, 3, -116, -128, 108, -110, 49, -66, 99, -42, 120, 20, -9, -87, -43, -54, 119, 70, 118, 82, -33, -55, -5, -51, -96, 63, -6, -114, 66, 127, -106, 34, 2, -94, 34, -18, -75, -44, 44, -104, 42, 37, 44, -94, 78, -126, -20, 70, 72, -30, 24, -88, 43, -108, -11, 75, 83, 111, 89, 22, 110, 111, -72, -16, -110, 91, 94, -57, -81, 11, -33, 89, -80, -116, 123, 126, -114, -25, 68, 86, 73, -35, 126, -12, -15, -12, -65, -60, -29, -104, 90, -46, -120, -109, 66, -102, 110, 33, -31, -99, -84, 64, 118, -36, 76, 114, -38, 90, -39, -97, 49, -93, -4, 47, 23, 109, -93, 87, -79, 7, 111, -116, 89, 119, -97, 27, -111, -115, -68, -14, -86, -24, -77, -96, 68, 127, -110, -97, 90, -20, -66, 11, 15, 58, -70, -90, 39, -34, 125, 88, 101, 109, 100, 62, 100, -125, -39, 118, -112, 22, -24, -70, 126, 27, -37, 67, 27, -19, 98, -11, 89, -96, -128, -24, 90, -70, 15, 1, 24, 12, -39, -3, -7, -66, -69, -34, -63, 21, -44, -46, -85, 60, 12, -87, -40, 103, 108, 115, -43, 78, -24, -82, 110, -24, 23, 72, 34, -90, -55, -69, 50, 35, 56, -84, 97, 116, 10, -94, 9, 94, -12, 52, 26, -127, 93, 114, 104, 74, 101, -67, 24, -51, -20, 7, 53, -125, -49, -40, -87, 25, 19, 91, -68, -53, -121, -99, -65, 17, -65, 72, -17, 52, -4, -118, 53, -38, 124, 29, -92, 98, 91, 60, -81, -57, -61, 101, -54, 19, -67, -13, -84, 80, -50, -24, -101, -42, 5, -37, 103, 68, -93, -41, -8, 32, -31, -83, 122, -35, 75, -98, -65, 38, 90, -17, 109, -98, -44, -73, 49, 17, 42, 93, -31, 120, -59, -4, -50, 74, 87, -74, 14, 123, 13, -121, 27, 110, -76, 21, -53, 127, 51, 11, 37, 13, 122, 18, 43, -50, 73, -36, 95, -13, -71, -64, -20, -2, 60, 58, -56, 20, 112, 87, 15, -3, 94, -86, -21, -110, 63, 55, -110, -14, -62, 55, 127, -68, -54, 43, 10, -109, -121, -23, 7, -63, 41, 115, 63, -27, 45, -120, 121, 30, 95, 8, -101, 61, 50, 7, 79, -15, -66, 97, 99, 0, 25, 99, 60, 99, 14, -58, 118, 21, 47, -3, 86, -40, -16, 22, 61, -98, 30, 55, 60, -3, -65, 87, -70, 114, -34, -119, -29, 28, 107, -57, -100, 4, -86, 88, -25, 56, -98, -35, -51, 77, 91, -92, -91, -53, 58, 99, -23, -40, 26, -91, 85, 89, 125, -113, 75, -37, -104, -81, 120, -125, -10, -108, 7, 32, 109, 110, -40, -117, -52, 37, 89, -89, 73, 126, -14, 3, 97, 92, 91, -5, -127, 48, -43, 126, 63, -96, -38, 88, -49, -46, 91, 69, -26, -29, -27, -45, -47, 61, -33, 29, -29, -72, 68, -84, -74, -73, 48, -104, -109, 11, 19, -108, -68, 104, -109, 123, -119, -19, 83, -40, 63, 47, -98, -91, -110, 3, -7, -29, -63, 88, -127, 36, -112, 69, 80, -58, 124, 0, -34, -113, -116, 114, -92, -56, 90, -73, -61, 99, 36, -105, -68, -29, 70, -38, 8, 88, 93, -127, -69, -98, 89, -68, 66, 105, -126, 19, -80, 126, -109, 14, -114, -97, 0, -78, -25, -37, -23, 43, -66, -115, 66, -6, -16, 8, 84, 120, -32, 50, 122, 27, 80, 83, 88, 19, 61, 90, -90, 109, 88, -71, -5, 102, -39, 124, -104, 64, -41, 1, -21, 21, 14, -83, -112, 126, 53, 100, 119, -107, 22, 113, 49, -25, 68, 9, 122, 1, -29, -96, -18, -69, -39, 106, -94, 50, 102, -70, -13, -67, 60, 94, 82, -54, -116, 98, -55, 65, 71, -64, 87, -35, -79, 8, 68, 117, -111, 62, -9, -12, 94, 101, 47, -72, 79, 81, 106, 53, -116, -35, 114, 72, -68, 69, -110, -56, 39, -37, -119, -18, 27, 96, 76, 76, -24, 16, 66, -7, -49, -71, 109, -83, -98, 29, -27, 110, -18, -48, 35, -6, 45, 22, -62, 105, -37, -43, -79, -126, 48, -69, -15, -52, -101, -67, -104, 4, 77, 90, 125, -100, -109, 107, -54, -78, 8, 47, -96, 118, 127, 67, -15, 45, -39, 51, 22, 52, -120, 72, 55, 57, -125, -88, -123, -98, -27, -99, 34, -78, 120, 32, -49, -117, 11, 25, -67, -109, -56, -35, -119, -56, -95, -6, 117, -6, -82, 11, -81, -74, -45, 102, 111, -42, -114, 116, -11, -13, -110, -105, 37, -118, 55, 116, -107, -62, 13, -45, -43, 86, 48, -33, -98, 81, 89, -109, -52, -121, 30, -5, -66, 114, -31, -83, -56, -17, -94, 61, 98, -76, 85, 7, -66, 12, -4, -45, 79, -119, 38, -92, 95, -41, 3, 125, -88, -35, -112, -12, -28, 47, 111, 34, 33, -48, 80, 105, 63, 114, 39, 33, -90, -4, -87, -28, -120, 37, 55, 87, 46, -34, 124, 14, 53, -1, 11, 93, 92, 28, -46, -63, -53, -63, 99, 108, 18, 51, 85, -47, 37, -4, 115, 75, 120, -100, -81, -127, 65, 103, 88, -17, -59, 84, 125, 122, -44, 9, 87, -80, -91, -87, -15, -16, -21, -43, -36, 125, -120, -79, -50, 46, 46, -63, -7, 38, -35, 41, 39, -98, 16, 0, 14, 85, -44, 11, 79, 40, -108, 38, 89, -71, 80, -54, 41, -69, 31, -123, -72, 40, -73, 6, -42, 101, 72, 79, 11, -91, -8, -77, -60, -120, 51, 82, 93, -121, -35, 44, 48, -14, -45, 9, 43, -93, 83, -43, -34, -13, -38, 22, -101, 17, -100, -15, -10, 100, -64, -126, -118, 57, -75, -50, 65, 104, -96, 31, 111, -3, -53, 31, 111, 30, -88, 27, 65, 124, 112, -97, -17, -54, 53, 10, 92, 82, 123, -46, 54, -69, -44, 64, 116, 9, -114, 54, -15, -82, -43, -31, 44, 32, -128, 27, -65, -87, -74, -128, -91, -90, -96, 20, -15, 85, -98, -51, 39, -103, 31, -34, -44, 116, -98, -55, -3, -83, 127, 111, -37, -44, -48, -121, 116, -48, 35, -77, -7, 89, -76, 30, -128, -44, -78, -15, -87, -48, 62, 81, -23, -35, -81, 62, -47, -51, -121, 79, -6, -122, 62, 86, -38, -114, 93, -50, -34, 0, 2, 88, -38, 54, -10, -38, -118, 41, 75, -77, 121, 9, -124, -29, 102, -77, -95, -72, 1, -88, -121, 123, -82, 69, 81, 8, 83, 47, 86, -79, -81, -40, -119, 9, -114, 0, 99, -104, -87, 46, -52, -94, -73, -48, 5, -98, 4, 38, -42, -123, 78, -35, -128, 124, -94, 82, 4, 117, 1, -37, -90, 48, 51, -80, -70, 66, 48, -99, 90, 89, 76, -90, 123, -125, -9, 1, -95, 123, -89, -9, -128, 118, 84, -128, 114, 118, 82, -9, 107, -45, 82, -110, -124, 5, -62, -66, -57, 114, -37, -94, 75, -89, -56, 70, -85, 63, -57, -52, 58, -17, 68, 58, -27, 24, 59, -41, 15, 13, 78, -6, 97, 32, 12, 101, -90, 78, -93, -19, 64, -2, 15, 11, 38, 88, -46, 81, 23, 25, -99, -46, -120, 97, -116, -19, -6, 71, 69, -119, -43, 19, 3, -74, -76, -112, -101, -38, 94, -66, 71, 31, 60, -41, -86, -30, -81, -4, -77, 70, -106, -47, -104, -98, -78, -91, 12, 44, 108, -47, 53, -63, 100, -71, -9, -104, -55, 18, -14, -89, 80, -70, 70, 13, 17, 113, 111, 64, -19, -93, 6, 3, -12, 31, 34, 38, 68, -82, -45, 48, -1, -120, 114, -29, -63, -23, -4, 10, 124, 110, 50, 76, -88, -8, -39, 57, -23, -55, -7, 87, -20, -128, -38, 96, 31, 124, 6, -29, -86, 89, -109, 41, 98, -123, -115, -93, -17, 9, 46, -21, -9, -32, -73, 32, 88, 17, -39, -62, 90, 83, -103, -58, 83, -13, -90, -14, -16, 44, 85, 26, 6, 104, -60, -24, 110, -47, 11, -35, 90, -71, 72, -47, 25, 127, 113, -14, 16, -53, 52, -22, -98, 77, 48, 113, -64, 86, -29, 48, 3, -72, -53, -119, -96, 15, -15, -114, 96, 124, -21, 58, -74, -77, -117, 79, -77, 125, -63, 67, -56, 117, -82, -26, 66, 94, -41, -125, 53, 58, 51, -72, 114, 126, -63, -110, 13, 50, -95, -19, 46, 12, -89, 100, 64, -77, 52, 115, -80, 117, 54, -8, 107, 100, 94, 45, 67, -75, 48, -8, 111, -28, 48, 97, -30, 113, 115, 112, 35, -108, -35, -47, 33, 5, -74, -31, 56, 106, -44, 104, 95, -118, -32, 74, 111, -66, -8, 50, -13, -88, -86, -30, 12, 90, -61, 111, 75, -74, 95, -18, -53, -68, 63, 108, 65, 117, -51, -7, 95, 33, -31, 63, 43, 65, 9, 26, 127, -127, -52, -14, -86, -10, 84, 54, -48, -105, 37, -101, -50, 4, 9, 25, 65, -55, 5, 2, -66, 82, 124, -98, -13, -35, 93, -98, -97, -26, 57, -98, -24, -123, 17, 18, -4, -27, -56, 76, -3, 110, 104, 75, -14, -15, -28, -77, 58, 105, 54, 121, 59, 50, -105, -82, -113, 116, -52, -82, -38, -123, -51, 66, -117, 94, -44, 7, -61, 29, -45, 64, 11, -69, 11, 125, 45, 111, -79, -25, 88, 103, -32, 19, 25, -9, 65, 40, -21, -114, 87, 70, -109, -92, 8, -98, -126, 93, 37, -59, -6, 121, -122, -123, -76, 17, -126, 97, 1, -77, -55, -39, -102, 41, 109, 51, -95, 46, -36, 12, 60, -77, -46, 80, -41, 91, 110, -39, 56, 20, 30, -78, 13, 36, -73, 65, -74, -71, 35, 55, -19, 108, -112, 7, 21, 125, -69, 54, 44, 23, -61, -24, 74, 21, -72, -95, -16, -89, -6, -88, 59, -104, -38, -56, 61, 17, -119, 115, 75, 44, 42, -72, 24, 58, 63, -82, 56, 122, 100, -28, 17, -89, 76, -37, 61, -123, -4, -83, -84, 118, -42, 103, -113, 48, -81, 76, -62, -72, 63, -115, 101, -23, -59, -3, -93, -124, 43, 91, 127, 16, -65, 16, 55, -116, 108, -12, -111, -24, 34, -67, -33, 120, -92, -18, 40, -45, -70, 106, 11, 121, 119, -16, -30, -68, 110, 5, -63, 25, -31, -64, -87, 32, 80, 97, 44, 60, -43, 61, -91, 119, 122, 4, 111, -98, 114, 24, -15, -84, 2, 125, -91, -6, -19, 7, 54, -37, -116, 119, 117, -19, -73, -98, -114, -120, 127, 58, 68, -43, -8, 105, -52, -14, -19, -68, 17, -33, 84, -126, 11, -42, 127, 48, 80, -19, -73, 7, 72, -60, -2, 61, 49, 54, 92, 63, 62, 91, -6, 2, -80, 114, -20, -3, -28, 89, 57, 117, -71, 13, 120, 68, 99, 119, -11, 52, -28, 44, -69, -83, 112, 57, 106, 34, -17, 70, -31, -83, 34, 91, 48, 82, 77, -100, -49, -78, 117, -120, -89, -82, 21, -97, 115, -7, -105, -24, -83, -5, -108, -24, 40, -123, -95, 19, 39, 17, -39, -120, 62, 123, 100, -18, 78, 49, 10, -99, 99, 0, -90, -117, 46, 59, -86, 33, -76, -63, -119, -31, 61, -98, 73, -27, -93, 107, 120, 74, -4, -46, 82, -70, -51, 54, 41, -101, -24, -77, -71, -53, 51, -33, -42, -30, -102, 1, -125, -49, 66, -115, 48, -1, -85, -6, 101, -50, -27, 93, -104, 97, -81, 106, -101, -3, 33, 68, 24, -119, 120, 81, -44, 43, -80, 43, -115, -53, -84, -111, 26, 110, -98, -54, -18, -55, 68, -45, 23, -87, -80, 47, -118, -32, 25, -90, 93, -70, 106, -11, -61, 98, -57, 24, 14, -9, -61, 27, 66, -17, 44, -36, -35, 74, 39, 75, -109, -21, -98, 42, 21, -49, -39, 31, 47, 115, 69, 12, -83, 48, -127, -15, 18, -56, -119, -96, 64, -52, 60, 2, 59, -24, 95, -104, -77, 6, 100, -58, 113, -126, 113, 6, -47, -54, -90, -128, -67, 107, 12, -21, 27, 14, 92, -82, 86, 101, -50, 22, -79, -118, -103, 108, -13, 120, -124, 38, -2, 104, 108, -17, 107, 93, 118, -68, -88, -100, -67, -27, -121, 73, 80, 35, -41, 44, 81, -82, 17, -97, 68, 66, -86, 93, 46, 29, 85, 51, -61, -45, 27, -81, 67, 6, -115, 57, 67, -75, 85, -128, 26, 92, 73, -21, -1, -95, -105, -48, -49, 41, -16, -109, -21, 26, 113, -102, -73, 70, 77, -6, -102, -24, 41, 93, 111, 54, 22, 50, 107, -21, 50, 6, -57, -5, 113, 71, 28, -120, -105, 107, 49, 7, 127, -99, -95, 112, -73, -40, 54, -124, 82, 80, -20, -4, 45, -37, -78, -61, -115, -98, 46, 63, 36, 118, -69, 21, 61, 87, 29, 84, 67, -49, -36, 66, -20, -3, 50, 35, 86, -24, 39, 40, -71, -109, -92, 102, -17, -41, -86, -4, -11, 88, -68, -103, 78, -9, 46, 11, -50, -53, -32, -111, 26, 60, 83, -122, -71, 5, 41, -113, 110, -48, 56, -89, -28, 92, -115, 83, -77, -73, -49, 40, -112, 11, 65, 94, -126, -17, -22, -47, 59, 74, -30, -43, 6, -74, -36, 63, 59, -123, 79, 41, -42, 7, 80, 58, -29, 94, 13, 23, -107, 92, -65, -91, -24, -127, -124, -22, -16, -18, 59, -85, -72, -98, 1, 62, -44, 93, -3, -113, 98, -52, 57, -72, 83, 9, 114, -73, -25, -1, 78, -3, -36, -115, 34, 68, -114, 38, -82, -1, -108, 106, 42, -52, -120, -85, -118, -36, -120, 8, -21, 107, 84, -92, -93, 40, 46, -106, 95, -107, 21, 45, 18, 113, 58, -75, 53, 73, 91, 100, -56, 112, 78, 114, -68, 86, -98, -57, -78, -90, 79, 29, -111, 35, 66, -75, -53, -16, -53, -86, 5, 96, 87, -104, 82, 18, -51, 7, -37, -88, -21, 35, -104, -71, 21, -43, -113, 51, 28, -63, 90, -21, 95, 107, -114, 33, -96, -38, -111, -21, 4, 22, -52, -36, 46, -98, 110, 123, 37, -55, -92, -111, 108, -68, -54, 1, 17, -38, -75, -83, 27, -113, 24, -6, 122, 39, -101, -101, -127, -84, 6, 5, 67, 82, 97, -15, 112, 79, -19, 22, -104, 17, 39, -124, 77, 113, 6, -33, -53, 59, 12, 103, 74, -91, -31, 68, 76, -3, 95, 77, 41, -26, -46, -20, -72, -76, 94, -87, -125, -53, 63, -100, 92, -26, -96, 41, -41, 38, -120, 35, -31, 21, 10, -85, 58, 107, 112, 6, -24, 79, -45, -110, -75, 37, -2, -18, 89, -36, 23, 93, 39, -42, 121, 3, 60, -103, -83, -109, 64, -75, 54, -95, 74, -64, -51, 4, -84, -67, -118, 20, -116, -35, 38, -62, -125, -91, 48, 92, 1, -57, 57, -87, 29, 50, 44, -39, 76, 89, -20, 12, -113, -93, 45, 89, -29, 122, -34, 15, -73, -24, -92, -60, 70, 74, 6, 73, 111, -74, 37, -15, -3, -33, 26, -102, -111, -58, -13, 93, -96, 95, -23, -81, -126, -105, -120, -26, -111, -26, 117, -55, 79, -103, 13, 21, 100, -109, -34, 83, -55, -125, -60, 70, -30, 94, 96, -12, -91, -45, -47, -59, -78, 59, -12, -75, 82, -4, 27, 99, 99, 16, -84, 50, 42, 57, -57, 14, 76, 37, -31, -107, 40, 38, 91, -117, 4, 59, -1, 41, -114, 80, 110, -63, 11, -30, -10, -35, 95, -111, -63, 66, 33, -19, -12, -53, -89, 59, 89, 115, -32, -69, -119, -120, 97, 100, -109, -27, 32, 18, -113, 46, -29, 125, 111, 110, -32, -27, -52, -65, -10, 13, -127, -104, 122, -11, -29, -95, -80, -67, -107, 16, -8, -98, 24, -39, -126, 44, 62, 34, -66, 77, -47, 33, 75, -64, 16, -85, 38, 92, -22, -100, -23, -21, -76, -29, 96, 24, 5, -112, 85, 26, 32, -51, 56, -72, 38, 58, 100, -28, -35, -93, -78, 46, 68, 125, 110, -44, -88, 20, -80, 18, 49, 25, 125, 101, 125, 93, -3, 2, 109, -46, -100, 13, 31, 84, 69, -59, 14, 42, 42, 107, 77, 92, 25, 17, 89, 8, 102, -127, -100, -106, 19, 77, 48, 16, 51, 45, -19, -80, -81, -38, 3, -53, 103, -94, -97, 44, -24, 45, -42, -110, 25, -93, 110, -78, 53, 71, 58, 27, 72, 87, 49, -37, 36, -31, 107, -41, -114, -40, 8, -67, 50, -117, 8, 25, -83, 39, -59, 21, -43, 28, 39, 110, 63, 21, -96, -12, -36, 91, -113, -92, 50, 65, -1, -42, -94, -22, 46, -79, 66, -74, -18, -12, -63, 119, -115, -18, 30, -45, -124, 115, 111, 43, 97, 46, -63, -126, -93, 29, 93, -78, 66, 15, 115, -63, 101, -106, 44, 19, -57, -18, 73, 53, 99, -118, 44, 112, -7, -53, -61, -3, -66, -78, -88, -96, 97, -23, -94, -124, -121, 127, -74, 73, 14, -86, -118, -13, -64, 54, -121, 7, -91, 80, -68, -120, 91, 105, 120, -44, -76, -68, 81, -14, -18, 121, 18, -49, -29, 52, -45, -22, 51, 10, -77, -63, 52, -67, 53, 116, 116, 60, -5, -103, 12, 55, -95, -25, 32, -103, 59, 84, -43, 12, -57, 68, 6, 89, -109, 105, 14, -25, -45, -63, 113, 6, 3, 37, 67, -72, 25, 55, 116, -108, 80, 0, 75, 113, 104, -20, -117, 35, -64, -32, -80, 7, -92, 54, -31, -72, 31, 111, 31, 114, -80, 16, -8, 51, -75, -69, 107, 78, 115, 95, 98, 67, -32, 45, 53, -56, -103, 64, 107, -38, -96, -101, 97, -59, 81, -62, -3, -16, -79, -100, -30, -30, 44, 90, -107, 97, -106, -127, 47, -119, 96, 17, 76, -64, -66, 1, 8, -40, -63, -12, 50, -30, 15, 19, 39, -31, 86, -92, 81, -121, -64, -76, -23, 108, -114, -1, 77, -92, 0, -4, -83, -32, -115, 122, 33, -53, -5, -87, 35, 61, 29, -43, -97, -83, 105, 70, 14, 63, 106, -33, 70, -86, 19, -80, -106, 34, 47, 99, 70, -81, -33, 116, 15, -20, 110, -80, 55, -23, -38, -37, -90, 119, 48, -59, -92, 25, -117, 50, -40, 117, -110, -97, -97, 37, -49, -75, -57, 126, -104, -114, -83, -9, -126, 60, 99, 112, 109, 27, -39, -57, 118, 0, -66, 38, 69, -29, -64, 81, -107, 24, 70, -89, 55, 102, 77, -122, -101, -108, -124, -76, -94, -79, 43, -92, 110, 15, -108, 91, -86, -18, -94, -96, 110, -32, 70, 51, 67, -122, 4, 89, 31, -53, -128, -42, -79, 77, -35, -52, 98, -31, 0, -124, 19, -84, -87, 1, 59, -67, -36, 101, 43, -2, -123, 25, 94, 75, -51, 34, 82, 81, -5, -15, -100, -5, 71, -51, -55, -92, 26, -85, 6, -102, -81, -103, -58, -40, 26, -127, 22, 118, 102, -63, -12, 107, 91, -46, 55, -88, 116, 9, 121, -17, 122, -106, 107, 65, -29, -76, 102, 125, -33, -20, -104, 14, 5, -34, 103, -97, -32, -3, -107, -58, 62, 9, -78, 25, 91, 105, 65, 80, -14, 59, -65, -20, 81, -86, -83, -76, -34, -109, -78, 61, -1, -54, -52, -124, 40, -77, -93, -120, 48, -72, -49, -18, 65, 1, -120, 29, -22, 73, -19, 92, 4, 44, -56, -43, 87, -11, 10, -75, 9, 60, 115, -120, -122, -65, -115, 46, -14, -80, 55, -94, -23, -122, 16, -86, 7, 24, 71, 113, -30, -76, 77, 102, 97, -107, -68, 56, 10, 70, 109, -109, 2, 96, -100, 8, -97, -87, -74, 17, -39, 109, 51, 66, 115, -60, 109, -6, 92, 52, -21, -66, 105, -72, -91, 74, -51, -31, 2, 88, -89, -17, 107, 41, -48, -121, -79, -17, -80, -25, -127, 10, -43, 52, -52, -56, 120, -71, 67, 85, 110, -82, -109, 87, -25, -72, 33, 52, 25, -93, 12, 64, 18, -8, -23, 98, -1, 26, -46, 48, -126, -45, -70, -41, -121, 6, 31, -128, 64, -30, 85, 46, 17, 104, 5, 120, -95, -90, 44, 58, -55, -71, -5, 91, 49, 100, 62, -80, -1, -112, 96, 1, -29, -102, 88, -22, 33, -9, -22, -31, 90, -65, -113, -21, -88, 20, -29, -55, 58, -113, -125, -125, -56, -2, 94, 121, -29, 28, -86, 98, 44, -118, -29, -113, -91, -69, -6, 70, 50, 100, -89, 12, -92, -74, 119, -52, 74, -38, 21, 4, -22, 24, 7, 50, -105, -27, 44, -6, -126, 86, -36, 46, 96, 63, 62, -123, 122, -72, 75, 44, -100, 114, -71, -64, -88, -80, 12, 114, 11, -95, -10, 117, 58, 125, 39, 81, -29, -45, -53, -27, -87, 39, -109, -118, -26, 81, -113, -32, -119, 91, -116, -90, 77, -59, -26, 118, -10, 115, 104, -127, -108, -33, 118, 78, -36, 29, 31, 63, 113, 106, -92, -102, 17, -72, -92, 119, -119, -76, -41, -109, -113, -28, -71, 92, 41, 31, 82, -97, 18, 59, -96, 39, -102, -106, -11, -10, 52, -107, -74, 37, 127, -38, 63, 17, 18, 100, 8, 28, -104, 96, 47, -89, -60, 104, -125, 109, 7, 86, -115, -102, 17, -83, 65, 43, -60, -74, -95, 120, -53, -41, 29, -53, 50, -36, 92, -60, -64, -28, 96, -40, -60, 15, -1, 8, -9, 3, -10, 127, -39, 3, -103, 106, 48, 90, 21, 116, -112, 54, 108, -36, -114, 9, 39, 64, 102, 3, -124, -90, 103, 101, -1, -84, -12, 126, 52, 108, 1, -86, 107, 90, 45, -124, 68, -34, 94, -39, -46, 110, -112, -65, -54, -98, 72, 113, 94, 46, -12, 98, 85, -36, 71, -44, 8, -68, -46, -68, -88, 84, -25, -109, 46, -108, -105, -13, -14, 117, 76, 69, 99, 92, -124, -82, 122, 76, -97, 88, -5, 20, 59, -48, 112, 2, 36, -8, 62, 118, 52, 102, 74, -101, 121, -7, -80, -112, 108, 34, -123, 56, -25, 105, 21, -21, -105, 15, -72, -74, -24, 51, 74, -93, -125, 58, 37, 39, -78, -28, 29, 103, -54, -24, -126, -60, 97, -78, -44, 77, 85, -38, 5, -68, -61, -102, 40, -38, 42, 96, 16, -110, 19, -37, -75, 22, -107, 90, -67, -56, -66, 90, -81, 9, -62, -79, 77, -93, -28, -95, 112, -71, -5, -10, -11, 62, 16, -99, -104, -70, 125, 41, -52, 16, -124, 1, -90, -103, -36, -29, -31, 26, -66, 16, -93, 0, 66, 112, 36, -90, -110, 20, -33, 13, -118, 84, -52, 27, 114, -28, 85, 111, -115, -94, 0, -111, 35, 38, -85, 127, -118, 12, 26, -56, -99, 61, 72, 95, 46, -20, -123, 64, -127, -28, -51, -117, -72, 25, 38, -86, 126, -4, -102, -117, 30, 26, -99, -63, -64, -56, -63, -54, 84, 91, 18, 113, 24, -37, 80, -58, 71, 85, -122, 72, -71, -44, 84, -14, 109, -6, 28, 107, 118, 54, 119, 20, -48, -108, 86, 17, -36, -105, 91, -80, 114, -18, -94, 10, 73, 114, 81, 16, 72, 87, -39, -127, -85, -83, -13, -103, 39, -112, -124, 30, 70, 123, -78, -105, -113, -120, 40, -21, -97, 3, 28, -111, 113, 62, 28, 58, 48, -19, -53, -8, -60, 36, -6, -16, 81, 109, 9, -8, 125, 13, -106, 68, 9, -55, 91, 24, -47, 3, -124, -15, -122, 32, 2, 120, -34, -98, 50, -114, 11, 125, 7, 80, 33, -127, -64, -14, 110, 73, 107, 108, -42, -127, 48, 95, -54, 11, -8, 28, -114, -4, -115, -108, -100, 15, -116, -6, 46, 63, 8, -71, 60, -113, -119, -34, -112, -55, 80, 127, -110, 59, 107, -23, 61, 27, -56, -121, -90, 64, 35, -76, -68, 48, -56, -40, -64, -43, 82, 110, -108, -37, -89, 80, -22, -79, -82, -5, -6, 127, -6, 13, 58, -27, 118, -9, -128, -66, -1, -90, 127, -94, -38, -69, 83, 34, 20, -109, 119, -26, -127, -117, 65, -88, 92, -84, -39, -118, 39, 84, -119, -95, -31, 68, 6, -41, -69, 6, 21, 58, 44, 20, 93, -122, 80, 48, 40, -28, 67, 32, 74, 68, 43, 12, 108, 7, 56, -58, 18, -33, -102, 27, 0, -5, -33, -122, 82, 27, 12, -25, -43, -72, 124, -78, -66, 76, 98, 102, -80, 37, 6, 122, -23, -78, 6, -42, 57, -66, 28, -53, 29, 54, 103, -99, -79, -58, -93, -125, 97, 47, -22, -73, 103, -26, -23, -91, -78, -52, -116, -30, 113, 18, -35, -37, 68, 99, 49, -2, -94, -51, 73, 63, -125, 48, 93, -76, 119, -128, -73, 88, 48, 33, -113, 23, -120, -7, 61, -70, 69, 73, 29, 54, -37, 122, -111, -96, 93, 66, 30, 127, -113, -25, 63, -110, -104, 28, -58, -113, 28, -3, 103, -52, -97, 119, 100, -89, -16, 33, -31, -75, -22, 126, 107, 69, 120, 125, 101, 86, 63, 3, 85, 79, 107, 20, 97, -125, -80, -88, -110, 77, 37, 121, -103, 68, 112, 125, 107, -32, 30, -51, 21, -120, -53, 1, 78, -60, -2, 51, -102, -67, -73, 111, -116, -94, 4, 110, -91, 52, -106, -73, 1, 59, -80, 27, 0, -95, 24, -21, 1, -73, 56, -105, -65, -124, 24, -115, -56, -106, 65, -30, -45, 120, -47, -32, -102, 85, -50, -65, 10, -28, -10, -117, -97, 38, 38, 31, 71, -65, -117, -55, -10, 67, -32, 53, 71, 120, 67, -113, -114, 4, -15, -31, -4, 67, 65, 22, 24, -113, 85, -94, -13, -53, -82, 19, 113, 84, -78, 57, -109, -67, -126, 9, -127, -30, -65, 72, -38, -126, 88, -24, 6, -55, 73, -126, -116, 11, 24, 37, 26, -19, 71, -114, 56, 117, 33, 41, 74, 83, -30, 93, -111, -28, -25, -110, 70, 38, 90, -96, 40, 50, 8, -82, 124, -46, -80, -120, 93, 72, 45, -9, -75, -11, 5, 109, -22, -90, 22, -76, 122, 121, -110, -117, -35, -7, -99, -92, -97, 119, -60, 71, 42, 77, 117, 38, -97, -91, 46, 124, 109, -36, -13, -94, 81, 121, -113, -69, -97, 37, -16, -103, 30, 2, -92, 124, 123, -63, -96, -102, -71, -28, 97, 99, -79, 86, 9, -48, 123, -73, -52, 104, 19, 64, -118, -28, 57, -103, 32, 88, 62, -112, 114, -35, 18, -106, -39, 13, -40, -7, 39, 17, 93, 8, -12, -113, -34, 125, -33, -39, -76, 44, -63, 72, -20, -53, -84, -91, -28, 76, 125, -94, 92, 111, -1, -18, -122, 88, 123, -34, -47, 34, 111, -81, -86, -29, -66, 8, -32, 29, 97, 20, -55, -94, -36, 53, -19, 9, 90, 81, -43, 88, 116, -78, 71, -13, 32, 77, -52, 28, -85, 29, -66, -102, 76, -23, -3, -118, 113, 93, 40, 83, -14, 113, 117, 78, 39, -29, -41, 1, -76, 45, -39, -88, 95, -95, 28, -1, 110, 104, -101, -102, 5, -38, -76, -46, 67, 50, -36, 52, 15, -124, 7, -127, 118, -3, 80, 29, 96, -89, -98, -108, 84, -8, -67, 51, 25, 89, -77, 7, 65, -50, 33, -58, 40, 86, 24, -21, 8, 117, -96, -105, 121, 39, -103, 111, -92, 105, 12, -124, -112, 43, -103, 101, -93, -42, 24, 60, -81, 75, -61, 112, -102, 101, -74, 66, 59, 79, -82, -61, 68, -50, -38, 61, 117, -13, 45, -102, -36, -71, -98, -19, 100, -73, -46, -121, 13, 106, 67, 60, 54, -121, 44, 80, 108, 99, 18, 39, 50, 64, 106, -10, -114, -60, -77, -124, 56, 96, -98, -108, -102, -68, 1, 126, -12, 83, -122, -127, 62, 73, 62, -12, 80, -22, -60, 60, -51, 86, -29, 127, 23, -51, -11, 37, 18, 41, 41, -54, 9, 71, -34, 35, -124, 96, 34, -8, 51, 40, -7, -15, -15, -73, 101, -62, 34, -87, 126, 111, -128, -30, 111, 23, 47, -28, -68, -63, -115, 102, 11, 23, 45, 106, -70, 49, 74, 92, -87, -3, 4, 35, 111, 118, 90, 84, -72, -4, 126, -74, -20, 126, 24, -37, 21, -56, 63, 81, 9, 77, 55, -107, -28, -27, 127, 30, -106, 73, -5, -64, -58, 127, 99, -75, 117, 61, -118, -83, -70, -120, -28, 38, -122, 124, -127, 27, -60, 64, -20, 78, 13, -92, 99, 113, 9, 98, 16, 31, 43, -117, 95, 113, -118, 66, -89, -128, 0, -79, -83, 58, -71, 17, -32, -65, 14, -31, 90, 82, -95, -58, 32, 47, -22, 3, 32, 115, -27, -80, 19, -112, -69, -14, -126, -58, -75, -87, -58, 53, -38, -13, -17, 19, -123, 79, 82, 19, -80, 44, -27, -47, 114, -122, -128, -35, 9, 33, -48, 111, 81, 99, 127, -115, -42, -127, -45, 11, -86, 25, -64, 4, -116, 47, -105, -111, -2, 105, 36, 46, 21, -118, 127, 8, -112, -128, 101, 25, 33, -75, 8, -14, -103, 8, -1, -17, 9, 82, 122, 52, -21, -70, -72, -8, 105, -48, 9, -25, -71, -82, -107, 79, -72, -108, -41, -56, -108, -68, 97, 53, -15, -22, -88, 10, 114, 39, 121, -5, -6, 115, -81, 101, -83, -24, -35, -106, 56, 103, -3, 113, -107, 18, 64, -51, 39, -105, 21, 59, -45, -10, -15, 69, 96, 25, -49, 82, -64, -55, -50, 58, -68, -3, 32, -22, 101, 125, 0, 29, 100, 126, 15, 121, 16, -49, -58, -73, -25, 91, 115, 58, -46, -28, -1, -78, 125, 79, -123, -67, -104, -45, 120, -44, 80, 24, 62, 54, 21, -65, -45, -6, -67, 98, -13, 77, -78, 58, -123, 25, 21, 120, -45, 103, -36, 83, -102, -39, 34, -97, 22, 58, -14, 14, -114, -62, -90, 77, 120, 60, -116, -52, -74, -55, -82, 41, -106, -32, -29, -101, 121, 121, -109, -51, 96, -17, -96, 122, 72, 66, -103, -33, -4, 11, 109, 10, 78, -108, -41, 70, 80, -29, -110, -122, 44, -63, 47, 67, 33, -109, 94, 27, -116, 114, 104, 108, -31, -120, 103, -86, 74, -128, 9, -58, 12, -10, 80, -38, 10, -88, -96, -38, 11, -77, -32, -72, -12, -112, 123, -107, -93, 89, 48, -81, 75, 24, -101, -83, 32, -126, -41, -22, -125, 96, 48, 15, -42, 1, 105, 97, 41, -119, -69, -76, -68, 28, -20, 48, 44, -25, 70, 79, -63, -10, 126, -116, -113, -103, -71, 47, -100, 16, -102, -97, -16, 74, 46, 71, -53, 23, 40, 116, 32, 99, -87, 93, -1, 21, 13, -85, 125, -45, 122, -66, 74, 120, -54, 89, -110, 4, 8, -82, -108, 34, -51, 5, -19, 123, -52, 56, 18, 116, 45, -78, 87, 86, -113, -41, -21, 29, 2, -24, 112, -3, 38, 58, -11, 113, 19, 7, -11, -100, 53, 9, 62, -126, -114, -85, 125, -38, 100, 15, -50, 17, 66, -90, -25, 81, -3, 82, -18, 127, -69, -33, -4, 97, -103, 114, 82, 45, -7, -57, 73, -81, 81, 7, -79, 95, 51, -81, -70, 23, 62, 8, -88, 0, 46, 15, -46, -85, -31, 64, -85, 28, -97, 39, -2, -71, 25, -48, 102, -109, 24, 47, -62, -23, -74, -13, -56, 105, 34, 2, 0, -31, -117, 40, 97, 57, -73, -77, 101, 25, 116, -112, -75, -109, 55, 51, -52, -47, -124, -78, -28, 28, 97, 38, -123, -104, -103, -51, -127, 60, 80, 2, -99, 91, -86, 126, 20, -30, -78, -7, 123, -90, 9, -80, -71, -63, 100, 6, 18, 104, 56, 118, 4, 26, 28, 9, 50, 53, 86, 51, -15, 38, -75, 14, 1, -32, 13, -106, 66, 63, 15, 61, 101, -103, 109, -98, -38, 81, 36, 108, 57, -35, 98, -67, 119, -2, 70, 41, -77, 29, -36, 37, -61, 18, -77, 69, 114, 64, 91, 52, -1, -22, -15, -28, 3, -34, 3, 93, -80, -89, 73, 105, 4, 43, -89, -5, -87, 109, -92, -35, 10, 1, -126, 78, -109, -75, 19, -123, 118, -18, 57, -11, 88, -86, 90, -36, 8, -35, -71, 56, 4, -125, 34, -119, 46, 73, 4, 88, 54, 41, -75, -63, -86, -73, -113, -67, -20, 34, -62, -30, -112, 123, 88, 104, -91, 50, -60, 45, -113, -2, -26, 19, 1, -120, 28, -81, 81, -95, -121, 7, 74, -68, 72, 116, -13, 87, -79, 96, -7, -13, -62, 9, -18, -102, -14, 19, 76, 54, -64, 91, -76, 38, -17, 53, 46, -117, 101, -1, -84, 108, -121, 118, -87, 79, 106, 28, 39, -101, -4, -96, 14, 63, 42, 124, 89, -100, 15, 38, 82, 80, 1, -121, -10, 112, 60, -91, 124, 33, 36, -88, 14, 43, -97, 55, -5, -119, -45, -94, -91, 80, -62, 51, 15, 108, 48, -24, -120, -65, -114, 91, -113, 16, 98, 6, 0, 30, 43, -4, -64, -49, 37, 78, 123, 68, 5, -10, 77, 88, 24, 114, 40, 90, 38, -73, 71, -42, 32, 79, 21, 46, 42, 37, -66, 12, -85, 63, -85, 86, -69, -21, -91, 96, -71, -96, 36, 62, 22, -14, 22, -82, -28, -65, -119, -118, -10, 80, -32, -106, 31, 118, 69, -54, 27, -125, 86, 70, 66, -127, 28, 126, -20, 65, 94, 37, 98, 3, -29, -8, 117, 122, 39, -39, -71, 48, -28, 47, 0, 68, 70, -97, 58, 11, -23, -43, 14, -64, -101, -47, -63, 55, -49, 46, -7, -83, -45, -37, 48, 55, 83, 37, 49, -6, 127, 106, -86, -29, 25, 42, -89, -33, 74, 98, 106, -77, -73, -7, -13, -45, 74, 53, -118, -103, -29, 3, -58, 54, 94, 119, -19, 50, 28, -98, -84, 27, -120, -41, 126, 34, -127, -90, -127, 75, -120, 108, 127, -65, -27, -14, 18, -81, -89, 29, -56, 10, -96, 14, -63, 127, 5, 46, 49, -94, 77, 93, 61, 85, -76, 60, -9, -74, 98, -7, -127, 106, -27, -128, -87, 74, -13, 60, 121, 26, -39, -63, -91, -7, 79, -26, -8, -43, -108, -87, -9, 97, -121, -76, 55, -69, 112, -82, -15, 82, 39, -13, 60, -116, -13, 102, 86, 102, 34, 79, 1, 123, -112, 38, -12, 96, -116, 109, -75, -96, -106, 44, -126, -99, 96, 57, -39, 81, 103, 74, 35, 15, -67, -32, 27, 49, -58, -14, 23, 104, -63, -104, 99, -46, 62, -41, -78, 74, -60, -25, 107, -37, -109, 109, -8, 115, 38, 81, 68, 13, 28, -24, -100, 89, 72, 56, 10, -114, -86, -94, 118, -21, -70, 89, 61, 121, -80, 111, 67, -11, -42, 46, 80, -23, 27, -56, -35, -63, -102, -95, 79, 54, 9, 107, 15, -47, 35, -102, -33, 77, -68, -43, -71, -10, -82, 118, -17, -33, 102, -77, 84, -68, 97, 36, 38, -3, 108, -125, 62, -122, -92, 13, 60, 46, -7, -52, 127, -100, -26, -33, 106, 34, 52, -93, -104, 99, -103, 8, -62, 127, 59, -106, -68, 28, 58, 98, -103, 38, 101, 88, 45, -119, -27, -23, 55, 94, 53, 55, 123, -101, -106, 101, 61, 74, -120, 86, 45, -95, -34, 111, -95, -103, -123, -35, 53, 63, -65, 79, -26, -92, 39, -109, -83, -116, -4, 101, 107, -78, 28, 102, -51, 50, 75, -117, -4, 83, 97, -86, 116, -65, -103, -107, -40, -97, -14, -115, 94, 49, 92, -60, 85, 3, -41, -125, 16, 84, 104, -5, -122, 4, -31, -45, -74, -84, -34, 50, 127, -65, 92, 115, -2, 118, -119, 86, -107, -5, 100, 115, -83, 64, -72, -126, -60, 15, -123, 84, -29, 109, -49, -23, -15, 48, 61, 39, 92, -101, -38, 91, -37, -74, 78, 89, -84, 87, 48, -63, -45, 20, -75, 0, -44, -19, 2, 24, 124, 8, -20, -32, -11, 59, 73, 103, -21, 6, 14, -57, 34, 104, -94, 125, -97, 113, 86, -53, 72, 6, 13, -101, -102, 66, 27, -17, -81, -98, -121, -85, 38, -12, 11, -101, -81, -43, -126, 27, 91, 17, 98, -3, -7, -123, -6, 24, 118, -47, 100, 62, 87, -15, 90, 114, -77, -11, -31, -30, 19, -24, 13, -71, 92, -103, -43, -116, -18, -41, 39, -55, 104, 9, 71, -30, 14, -63, 122, 4, 18, 94, -61, -22, -49, -99, -36, 2, 18, 61, 100, -90, -91, -14, -33, -126, 11, 52, -114, 121, -116, 53, -62, 116, -66, -119, -42, 77, -53, -47, -47, 93, -81, 20, -57, -1, 49, 35, -127, -60, -32, 102, -22, 6, -40, 73, 8, 99, -2, 22, 92, 10, -53, -98, -2, 9, -88, 85, -42, -13, -90, 40, -48, -43, -68, 24, 84, 110, -69, 86, -78, 28, 60, 28, -94, -108, -27, 42, 119, 99, -64, 83, -19, 11, 113, 108, -108, -103, 65, -21, 12, 103, -109, 93, -68, -49, -11, -111, -67, 48, 103, -17, -52, 35, -117, -18, 55, -15, -104, 46, -44, -40, 1, 66, 99, -14, 46, 120, 12, -17, -29, -104, -42, -10, 117, 18, 69, -22, 35, -125, -101, 10, -14, -25, -83, -2, 86, 100, 111, 110, 18, -61, -57, -109, -123, -86, 6, 51, -94, -110, -94, 5, -86, -8, 123, -96, -117, 65, 10, 46, 68, 37, -71, -74, -115, -26, 52, 99, -53, 35, 81, 93, 103, -104, 113, 108, -61, -9, 32, -27, 9, 66, 107, 51, -69, 102, 83, -58, 39, -34, 116, -21, -125, -83, 34, -112, 20, -42, 115, 95, 122, 69, 60, 97, 93, 45, 77, -96, -92, -19, 6, 45, -80, -15, -31, -21, -41, -76, 49, 127, 18, 37, -22, 22, 83, -116, 38, -25, -29, 26, -58, -35, -33, -126, -66, -68, 48, -117, -35, 84, -7, 99, 2, 41, -44, 99, -108, 43, -105, 69, 42, 42, -22, -107, -64, -67, -95, 102, 36, 4, 0, 106, 97, 95, 109, -97, -100, 29, -85, -7, -15, 36, -36, 115, -51, 48, 86, -31, -37, 110, -90, -122, 24, 16, -101, 88, 78, -68, 62, -14, 65, -65, -35, 34, -98, -54, 66, -70, 103, 109, 51, -40, 17, -113, -52, 94, 63, -94, -65, -101, -112, -27, -95, 40, 117, -68, 0, 67, -8, -65, -74, -71, -2, 19, 92, 28, 93, 30, 87, 68, 11, 10, -100, -100, 26, -24, 122, -39, 11, -71, -12, 27, 30, 21, -60, 19, 81, 68, -41, -54, -125, 13, 3, 1, -96, -33, -98, 125, 125, 117, 65, 8, -1, 93, 36, -103, -58, 30, -13, 81, 87, 103, -20, -11, -3, 48, -119, -50, -11, -32, 24, -8, 109, -100, 122, -115, -5, -104, -118, -7, -115, 75, -127, 12, 40, 38, 38, 110, -60, -103, 63, -100, -128, -84, 17, -3, 92, 26, 76, -47, 122, -28, 74, 103, 0, 68, 116, 124, 92, 126, -11, 105, 73, -10, -11, -14, -100, -101, -32, -31, -76, -96, -3, -75, -52, -114, 50, -88, 41, -2, -6, 35, 99, -60, 11, -29, -120, -1, -33, 100, -2, 84, 77, -57, -53, -62, 57, -25, -34, -102, 72, 18, -70, -59, 71, 6, -44, -6, 46, 125, 120, -88, 32, 91, -20, -85, -65, -12, 43, 30, -40, -87, -13, -91, -16, 62, -24, -86, -91, 70, -60, 110, -40, -2, -77, -96, -124, 7, 26, 50, 4, 18, 91, -91, -18, -57, -48, 45, 60, 123, -53, -108, -92, 62, -70, 21, -4, 34, 63, 34, -24, -125, 16, 64, 1, 67, 96, 5, -53, -6, -73, 79, -115, -110, 116, -5, -38, -59, -88, -106, -64, -13, -86, -27, -78, -28, 122, 46, -122, 57, -48, -18, 60, 96, -81, -67, 36, -113, 66, 111, 10, 121, 62, 23, -116, 51, -110, -26, 120, -70, -4, -72, 45, 38, 29, 95, -117, 23, 14, -111, -48, 94, 0, -116, 63, 47, -55, -29, 62, -117, -46, -56, -123, -112, 95, -111, 67, 113, -9, 59, -85, 115, 116, 89, 25, 17, 56, 36, -87, -58, 54, -7, -91, -74, 6, 100, 101, 79, -57, 35, 91, 25, 108, 96, 41, 75, 113, -19, 61, -24, -88, 104, -37, -100, 65, 116, 46, -6, 25, 87, 64, -49, -48, 101, 5, 86, 73, -22, 38, -112, -115, 1, 41, 121, -31, -45, 69, -46, 64, 2, 58, 104, -22, -107, -123, -84, -119, 51, 38, 34, 10, -26, 113, 90, -52, -10, 49, -107, 96, -41, -90, 110, 88, 79, 103, -71, -94, 44, 11, 98, -82, -59, 75, 25, -38, 80, 69, -29, 3, -21, -122, -115, 81, 119, 103, -99, -18, 24, -77, -50, 111, -39, -68, 71, -88, -92, -128, -53, 80, 11, -83, 127, 80, 120, 24, -86, 72, -35, 14, -53, 72, 20, -40, 25, 11, -64, 55, 121, 88, 106, -56, 72, -61, 4, 15, -21, 40, 16, 54, -7, -101, 100, -8, 108, 92, -112, -106, 37, -19, 36, 112, -75, -72, -55, 78, 68, 9, 5, 61, -31, -17, -123, -87, 50, 10, 57, -98, -78, -55, 84, 43, -28, 56, -93, -48, 21, -77, -25, -70, 32, -117, -86, 85, -60, -13, 36, -120, 124, -87, 69, -34, 25, 75, 7, -53, -43, -64, -23, 7, 9, -66, -77, 110, 118, -42, -66, 11, 10, 37, 69, -86, 49, 112, -128, 117, -29, 36, 125, -32, 77, 66, 62, -26, 13, -59, 50, 98, 6, -101, -22, -113, -39, 29, 125, -48, 115, -68, 91, -3, 97, 33, 40, 18, 17, 40, 7, 116, -52, 4, -44, -103, -57, -110, 0, 84, -40, -78, 55, 94, -51, -95, 109, 39, 62, 107, 119, 49, -89, 82, -81, -120, -13, 87, 27, -124, -1, -94, 121, 75, 39, -51, 100, 110, -32, -28, 66, 56, 22, -7, 22, 100, 26, 3, 11, -40, -18, 2, -118, 21, -44, -71, 30, 72, -112, -71, 76, 15, -37, 69, -38, -126, -109, -66, 112, -13, 35, 51, -85, -71, -84, 65, -99, 71, -60, 40, -97, 51, -86, -87, -56, -1, -30, 102, -57, -14, -97, -109, -127, -5, 89, -37, -3, 108, 26, -18, -33, -67, -95, 10, -10, -51, -53, 20, -108, 15, -68, -76, -62, -25, -35, 11, 102, 64, -15, -83, -78, 17, -64, -76, -116, -103, 15, 9, -123, -87, 119, -28, -26, -104, 110, 93, -26, -71, -15, -6, 73, 45, 46, -117, -108, -116, 22, 122, 76, -120, -89, 126, 25, -24, -78, 37, 1, 66, -82, 7, 107, -90, 107, -46, -66, 90, -81, 36, -109, 32, -97, 92, -51, 77, 104, -30, 89, -2, -36, 37, 6, 4, 36, -97, 108, 86, 68, -19, 24, 115, 116, 4, -103, 96, 86, -41, 58, -123, 124, 77, 37, -101, 42, 114, 104, 18, -44, 66, -112, 49, -25, 23, -75, -117, 54, -95, 98, -5, 14, -6, -18, 3, 126, 7, -29, 84, 94, -99, 89, 90, 106, -2, 117, 20, -15, 94, -90, 69, 32, -73, -10, -121, 78, 43, -109, 4, 76, 117, 127, -37, -17, -19, 94, -18, 116, -63, -62, 83, -34, -100, 45, -56, 26, 35, 93, -117, 1, -125, 81, -95, -70, -57, -88, -120, 115, -69, 13, 63, -80, 12, -102, 32, 122, 120, -114, 110, -71, -48, 65, 23, -20, -17, 96, -121, -110, 61, -110, 19, 64, 99, 52, 123, -85, 92, -125, -98, -104, 16, 93, -56, -99, 120, 104, -105, 112, 118, -123, -86, -57, 71, 65, 51, -74, 33, 58, -56, -34, 77, 91, -97, 48, 15, -102, 91, -21, -99, 121, 3, 46, 87, 76, 75, 79, 52, 98, 63, 43, 103, 105, 114, 46, 43, 37, 100, -52, -32, -84, 43, -83, -121, 74, 93, 22, 100, 57, -126, -127, 50, 5, 47, 9, -47, -6, -40, -122, -36, -104, 49, -60, -127, 35, 114, 44, -56, 87, 121, 40, -125, 36, 85, -117, -18, 51, 33, -46, -20, 35, -45, -98, -87, -125, 40, -6, -3, -128, 0, 90, -104, -79, -98, -102, 84, -112, 70, -99, 103, 63, 69, 107, -29, 27, 118, 81, -50, 23, -93, 58, -69, -9, 88, -28, -6, 0, 94, 119, 1, -33, 81, 25, 16, 111, 51, -27, -128, -6, 2, 103, -71, -57, 82, 29, 98, 72, -18, -80, -32, 18, 106, 27, -119, 67, 127, 3, -61, 93, -6, 68, -68, -52, -34, 77, -69, -111, -78, -69, 11, 52, -93, 69, 123, 117, -30, 94, 62, 80, -114, -98, -30, 121, 57, -21, 60, 56, 110, 127, 21, -23, 68, 82, 53, -94, 31, 112, -77, 81, -84, 63, 5, -49, 4, 0, -60, 102, -34, -126, 54, -19, -96, -103, -26, 89, 4, -94, 17, -13, -95, -89, 92, 101, 121, 17, -121, 24, 1, -69, -23, 45, 122, 110, 124, -2, -18, -63, -28, 77, -61, -102, -70, -28, -77, 32, -67, 56, 66, 79, -85, 99, 118, -121, 73, 111, 24, 80, 7, -103, -117, 112, 71, -123, 94, 67, 3, -52, -124, 103, -103, -56, -126, -45, 44, -75, 115, 105, 109, 53, 56, -104, 25, 46, -97, -30, 29, 55, -78, -92, 81, -66, -108, 24, -61, 114, -37, 71, -65, -32, 46, -40, 40, 48, 44, -44, 102, 31, -67, 83, -43, 118, 108, 110, 36, -117, -48, -62, 67, 2, -26, 20, 64, -5, -84, -124, -19, 7, 75, 44, 103, -7, -123, 15, -86, 49, 99, -112, -48, -95, 99, 37, -105, 79, 19, 59, 91, 99, 125, 30, -26, -28, -78, -90, 95, -34, -86, -52, 101, 117, 121, 77, -17, 126, -36, 25, 47, -64, 41, 127, -31, 12, 37, -8, -36, -72, -77, -73, -100, -79, 85, 2, 21, -121, 40, -12, -27, 83, 64, -54, 72, 57, -105, -73, 55, -12, 80, -26, 52, -7, -26, -107, -122, -117, 13, -30, -61, 64, 25, -33, 113, -18, 97, 6, -11, 10, 122, 90, -35, 59, -92, -91, -12, -68, -35, -84, 48, -83, 18, -28, 39, 120, -7, 45, -125, -122, -113, -57, 70, 40, 38, 56, -106, 8, -66, 11, -110, -71, -27, -17, 116, 9, 20, -24, 69, 113, 20, -11, -97, -89, 89, 70, -97, -46, -13, -93, -40, 2, -22, -97, -86, -112, 87, -64, 24, -107, 75, 42, -50, -80, -103, -62, 57, 46, 43, -1, 31, -65, 116, 62, -26, 78, 4, 6, -96, 119, 41, -7, -7, -109, 24, 35, -93, -17, 99, 60, 4, 46, -26, 83, 94, 0, -107, 24, -82, 64, -105, 77, -128, -117, 12, -26, 89, -112, 108, 122, -120, 21, -13, 1, 40, -117, -91, 76, -6, -120, 8, 126, 55, 110, 81, 21, -18, 103, -83, 28, 39, -60, -22, 39, -48, 118, -114, -87, -122, 122, -93, -114, 16, 22, 16, -72, 33, 53, -124, -101, 61, 12, -102, -12, -5, 107, -118, 105, 82, -73, 6, -6, -4, 112, -95, 76, 102, -81, 117, 108, -86, -103, 123, 58, 47, 11, 114, -47, -64, 119, -20, 125, 3, 6, -14, 126, -14, -4, 104, -60, 51, -18, 62, -81, -34, 96, 123, -60, -113, 113, -80, -71, -118, -85, 115, 57, 54, 102, -118, 118, 93, -9, 116, -32, 125, -26, -33, -17, 98, -57, 52, 21, 53, -14, 69, -109, -46, 64, -41, -30, 49, 7, 27, 59, 51, 15, -11, -23, -11, -1, -32, -46, 118, -44, 50, 116, 58, -111, -29, 28, -40, -105, -79, -115, 10, 118, -96, 92, 55, -9, -66, -24, 127, 90, -92, 50, -23, 25, -101, 94, -104, -5, -80, -113, 79, 98, -125, 9, 116, -26, -91, -52, -2, -41, -38, -120, -51, -6, 100, -124, 114, -93, -19, 113, 125, 17, 35, -26, -86, 62, -60, -62, -70, -12, -47, -119, -42, -44, 19, -54, 59, 56, 23, -71, -113, 113, -63, -35, -21, -91, -31, -35, -56, 78, -50, -59, -33, 113, 43, 9, 48, 111, 76, 106, -29, -99, 115, 58, -14, 6, -124, -83, -65, 27, -26, -50, 12, 39, 43, 120, 76, -115, -43, -107, 91, 36, -38, -69, 21, -122, 68, -59, 117, 16, -81, -39, 46, -93, -109, -96, 41, -105, -51, 104, 51, 51, -73, -65, -38, 98, -73, -90, 111, 13, -69, 75, -79, 22, -122, 70, 28, 74, -116, 17, -37, -69, 106, -119, -34, 125, -87, -120, -107, -10, 112, 72, -87, -89, -121, 3, -118, -65, 41, 121, 76, 101, 68, 125, -5, 74, 67, -105, 21, 79, 40, 112, -117, 19, 121, -23, 16, -94, -15, 37, 24, -30, -19, 65, 9, -11, -60, 19, 52, 109, 13, 0, 82, -47, -3, -51, -100, -64, -28, 49, -112, -115, 33, -101, 32, 26, 4, -80, 60, 118, 86, -44, -40, -61, -107, 97, 56, -39, -11, -20, -58, -126, 108, -103, -45, -23, -26, -17, 42, 75, -96, 58, 88, 65, 85, -8, -37, -39, 40, -105, -49, -2, -21, 39, 66, 0, 9, -6, 89, 126, 103, -96, -128, 83, -71, -45, -67, 31, 67, 103, -22, 99, 33, -62, 37, -10, 58, -128, 79, -29, -104, -97, 97, 3, 70, 35, -124, -49, -98, 93, -51, -123, 125, -51, 88, -74, 33, -107, 86, -28, 124, -64, -57, 29, 3, 108, -109, -67, 109, 99, 32, -123, -126, 2, 8, 72, -91, 12, -104, -61, -22, -27, -56, -25, 51, -95, 30, -44, -74, -12, 56, -77, 52, 127, 80, -73, 108, 100, -11, 89, 71, -107, 94, 73, 23, -26, 17, 61, 115, 41, -128, -35, -113, -55, 68, 66, -22, -30, -106, 32, 86, 78, 83, 11, 77, 36, 66, 57, 8, -73, 18, -49, -51, -16, -104, 100, 87, 41, 33, 74, -45, 34, -89, -30, 107, 107, -92, -43, -50, -70, 117, -92, -120, 73, 47, 85, -19, -14, 15, 117, 41, -95, -60, 118, 18, -36, 91, -23, -123, -4, -77, -40, -98, -38, 58, -119, -59, 94, -34, 19, -104, -44, 56, -96, -99, -25, 118, 10, 89, 5, -1, 3, 38, 67, -7, -72, -97, -44, 33, -92, 81, 84, -3, 111, -82, -73, 121, -12, -106, -41, -121, -82, 43, 63, -49, 72, -89, -59, -46, -128, 74, 81, 3, -16, 20, 125, 41, 51, -47, -54, 88, -94, -97, -43, -110, -51, 12, -117, 65, 34, -30, 73, 81, -114, 8, -96, 86, 47, -27, -87, 48, -81, 122, -77, 31, 15, -80, -56, -62, 2, 19, -102, 36, 50, -17, 54, 127, 124, 65, 65, 30, -92, 10, -17, -78, -110, 15, -120, 66, 116, -79, -14, -93, -84, 37, 67, 59, 86, -117, 125, -40, 30, -104, 124, -48, 7, 51, -48, 3, -12, -111, -94, 24, 27, 17, 74, 45, -95, 83, -17, -107, -124, 97, -71, -80, 7, 124, 107, -35, -121, 105, 53, 38, -127, 49, 118, 8, -28, -58, -116, 89, -41, -82, -15, 114, 63, -68, 32, 96, -113, -113, 118, -109, 113, -81, -60, -8, -85, -81, 85, -78, -104, 10, 88, -103, -69, 79, 34, 32, -107, 46, -7, -19, 92, 106, -33, 27, -90, 127, -4, -75, -113, -14, -55, -128, 33, 13, -8, 76, 60, -51, 126, 85, 87, 87, 110, -110, 38, 16, 50, 59, -66, -85, -88, -102, -106, 8, 54, -68, 7, -78, -14, 22, 36, 59, 22, -59, -56, -114, -111, -124, -37, -113, 89, -78, 102, 72, -59, 12, -40, 119, -56, 23, -93, -16, 49, -71, 120, -25, -11, 0, 25, 103, -106, -67, 34, 45, 2, 106, 59, 19, 111, -105, 35, 72, -55, 9, 16, 14, -106, 105, 6, -34, 0, 41, 78, -79, 98, 71, 25, -41, -57, -78, -65, -35, -16, 97, -118, 114, 76, 70, 6, 59, 93, -87, 3, -90, 50, -108, 53, 72, 125, -69, -90, -3, 100, 117, 46, 70, 60, -57, -99, -125, -6, -36, -32, 106, -66, -21, 92, -118, -79, -30, 69, -114, 11, -56, -76, -66, -36, 105, -122, -39, -92, -83, 86, -120, -94, 5, 78, 94, 76, 108, 97, -58, -56, -63, -80, 6, 44, -115, 16, 93, -17, -43, 107, 123, 30, -96, -71, 122, -119, -65, -44, -82, -20, -86, -74, 14, 47, -123, -20, -4, 113, -51, 66, -71, 15, 115, 64, -69, -128, -48, -103, -17, 38, -124, -22, -60, -92, 35, -66, -82, 99, 18, -36, -49, 61, 18, 94, -20, 23, -54, 104, 8, 24, 43, 66, -89, 30, 2, -30, 30, 82, -5, -115, -8, 0, -8, 60, 36, -101, 123, 82, 126, 13, -82, -50, -54, 65, -84, 55, -40, -10, 31, 97, -114, -54, 35, -75, 104, -91, 24, 6, 119, -109, 20, -16, 19, -116, -84, -72, -89, -89, -118, -90, 53, -71, -12, 127, 122, 32, 54, -46, -106, -42, -77, -91, 32, 86, -38, 9, 123, 114, -113, 115, -122, 35, -29, 25, 47, 15, 81, 87, 55, 92, 125, -20, -107, -15, -21, -113, -111, -94, -31, -89, -8, 21, -52, -104, -21, 39, 33, -25, 25, 49, -38, 31, -44, 61, -71, -124, -52, -118, 91, -125, 102, 88, -17, 123, -55, 91, -118, -38, 125, -20, 1, -11, -127, 78, 13, -20, -11, -81, 83, -114, 96, -83, 46, -76, 106, 103, -72, -73, 113, -109, -70, 88, 107, 42, 83, -76, 5, 94, 14, 2, -54, -112, 119, -53, 94, 4, 55, -45, 51, 11, -31, 19, 56, -113, 72, 35, 118, -128, 90, 104, -108, -108, 64, 127, 62, 19, -76, -61, -15, 66, 69, 59, 82, 60, -122, 48, -63, 62, -125, 116, -55, -27, 8, -127, -12, -48, 36, -21, -48, -2, -45, -28, 19, -109, -28, -47, 38, 24, 21, -104, -38, -38, 83, -83, -105, 90, 93, -40, 24, 97, -52, 97, -58, 84, 98, 58, -92, 7, -91, -11, -123, -8, 89, 24, 11, -67, 106, -78, 85, -1, -54, -80, 89, -99, -35, 112, 119, -70, -56, 15, -101, 21, -16, -31, -23, -45, -100, 14, 90, -63, -125, 95, 58, 92, -8, -59, -102, -30, -9, 111, 97, 65, -97, 58, 95, -4, 43, 86, 55, 115, -26, 82, 8, 86, -76, 114, -87, -48, 0, -125, 17, 3, 99, -53, -33, -37, 17, -7, 61, -120, -23, 30, 74, 8, -40, 41, -123, -125, -1, 60, 119, 101, 14, -1, 60, 66, -15, 101, -110, 113, 105, 36, -12, 76, 111, 84, -89, 0, -51, 100, 9, 54, 2, -45, -65, 90, 124, -60, 94, -5, -128, 85, -31, 14, -44, -99, -47, 70, -126, -29, 55, 107, -121, -84, 55, 119, -128, 94, -9, -51, 66, -128, -124, -60, -45, -61, -97, -49, 7, 125, 75, 7, 82, -84, -107, -90, -55, -26, 108, -53, 74, 36, -73, 81, 80, 110, 72, 80, 77, -64, -99, 15, -64, -95, 84, 20, -28, 115, 99, 107, 112, 46, -14, 66, 90, 8, 104, -93, 110, 85, -17, 56, -7, 38, 10, -55, 20, -46, -103, -31, 18, -74, 113, 83, -40, 69, -25, 60, 56, -54, 40, 40, 121, -102, -22, 83, 34, -46, 119, 17, -89, -26, -55, 32, -116, 83, 105, 32, -90, -126, -126, 56, -71, 115, 11, 17, 56, 114, -51, -16, -67, 117, -104, -74, -112, 2, -119, 50, 84, -128, -61, 124, -26, 13, 28, -14, -32, 6, -109, 6, 8, -107, -65, 65, -120, 74, -46, 64, 61, 32, -80, 122, 21, -56, -80, 37, 74, -71, -40, 30, -70, 27, 26, 32, -88, -73, -109, 9, 61, -90, -113, -59, -69, -50, -121, -61, -103, -39, -125, 86, 121, -77, 80, 15, -5, -128, -76, -59, -71, 12, 99, -13, -88, -2, -108, -48, 53, -89, 89, -14, -51, 105, 55, 8, -73, 62, 75, -48, -104, 78, -90, -111, -127, 118, 32, -4, 118, 85, 65, -80, -31, 36, 35, 9, -94, 55, 90, 87, 94, 51, -55, -85, 28, -127, 51, 84, 63, -2, -92, 87, -52, -53, 105, -51, -63, 9, 73, -72, -34, 10, -24, 64, -81, -117, -55, -47, 67, -93, -87, 33, 87, -14, 77, -13, -13, 0, -57, -77, 127, -20, -118, -53, 55, 115, 25, 120, -3, -30, -80, 91, 109, 24, 27, -100, 36, 101, -19, -25, -120, 22, -120, 95, -119, 85, -45, -4, -42, 26, 47, -43, -122, 58, 32, 61, 45, -71, 54, -86, 28, 102, -122, 9, -1, 33, 37, -93, 6, -110, 10, 15, 41, 18, -18, 50, -24, 65, -82, 62, -36, 94, -109, -30, 24, 51, -96, -59, 109, 86, -16, 9, 60, -10, -110, -69, -105, 55, -34, 30, 73, 104, -83, -14, -5, 27, -92, 99, -35, -45, 33, 57, -79, 52, -101, 73, -25, -69, -114, -44, -111, -2, 93, 78, 116, 111, -119, -116, 38, -24, 42, -16, -48, 87, 98, 75, -14, -121, 46, 79, -38, -49, 8, 11, -125, 36, -44, -21, 95, -30, 63, 113, 97, 29, 63, 85, 12, 72, 97, -77, -80, 11, 35, 1, -30, 5, -52, 85, 12, 123, 36, 102, -54, -83, -15, -50, 81, 69, 57, 48, -88, -8, 33, -119, -107, -32, 94, 34, -87, 64, 85, -39, -53, -8, 90, 46, 125, -89, 3, 10, -94, -89, -16, -20, -44, 98, 58, -91, 39, -13, 86, 79, 108, -9, 88, -127, 88, 55, 35, -127, -9, -8, -38, 66, 112, -75, -16, 110, -36, 115, -8, -2, -101, 104, 106, -17, 74, 37, 21, -14, -104, -21, -63, -124, 98, -102, -122, 58, 81, 41, 59, -56, -94, -106, -118, -110, -53, -5, -128, 39, -18, -8, -91, 9, -31, -113, 121, -85, 52, 14, 29, 77, 121, 95, 81, 91, 121, 87, 22, 74, 1, -47, -110, 35, -25, -100, 53, 50, 23, 54, -39, -122, -82, -2, 15, 15, 14, 8, 59, -62, -106, -40, -113, -113, -73, 97, 107, -80, 56, 1, 122, -71, 82, -116, 92, -70, -87, 18, 108, 64, -56, -58, 70, -10, 68, -42, -122, -46, 94, 65, 21, 117, -103, 36, -124, -47, 5, 111, 1, -66, -16, -4, -9, -61, 8, -44, -3, 49, 102, -23, -14, -82, 47, -72, 36, -12, 14, 42, 70, -19, -21, -37, -30, 5, -128, -26, 86, 5, -42, -41, 67, 70, 83, -69, -119, -36, 15, 6, -115, -11, 112, -1, 35, 31, 56, -57, -109, -58, 114, 90, 51, -35, -75, -107, 98, -75, -4, 56, 59, 82, -112, -2, 24, 99, 57, 34, -65, -56, -88, -51, 61, -104, 76, -32, 56, 4, 40, 75, 75, 26, 37, -2, 119, 91, 20, 90, -112, -112, 18, 75, 98, 34, -54, -6, 6, -125, -100, 69, -52, -59, -110, -119, -35, 95, -22, -107, -29, -110, 97, -82, 44, 6, 45, 35, -31, -63, -3, -14, -47, -112, -67, -77, 50, 7, 45, -72, 11, 74, 126, 87, -113, -112, 96, -20, 111, -54, 2, -45, -36, -29, 1, -120, 105, -82, 44, -53, -17, -87, 61, 64, -71, 122, 115, 108, 2, 33, -92, -115, -21, -94, 100, -6, -77, 68, 102, -94, -113, -24, -11, -21, 75, 119, -12, 53, -91, -96, -128, 21, -55, 61, -43, 3, 55, -55, -17, -71, 106, 19, -58, -43, 54, -86, 79, 105, 111, 53, -117, 126, -98, 1, -23, 105, -8, 93, 30, 29, 125, 30, -78, -57, -37, 8, 74, -109, 81, -71, -52, 59, 76, 19, -112, 2, 61, 95, -21, 44, 20, -9, 42, 50, 120, -108, 28, -16, 113, -70, -115, 111, 89, -64, -74, -76, 72, -128, -57, 25, -71, 20, -44, -123, -89, -28, 8, 100, -61, 115, 17, 87, -22, -69, 10, -30, -49, -90, 82, -63, -32, 96, -80, -71, -96, -26, -18, 104, -26, 53, 1, 31, -55, 85, 36, -16, -71, -84, -43, -4, -96, 102, -45, 10, -95, 93, 109, -15, -125, 63, 50, -28, 31, 98, 29, 63, -56, -117, 39, 46, 65, -88, -51, -118, 125, 113, -5, -74, -98, 80, 50, -66, 54, -122, 72, 87, 99, 53, -56, 103, -11, 122, -53, -108, 92, 104, 84, -92, 116, -5, 82, 53, 36, -97, 63, 33, -111, -70, 88, -81, -118, 10, -19, 64, 16, -75, 24, -12, 107, 96, -37, -32, 91, 38, -12, 55, 14, -56, 92, 2, 68, 46, -73, -24, 78, 119, -119, 95, -79, 97, -114, -68, -20, -5, 124, 124, 48, 20, -16, 27, -11, 75, 123, -48, -15, -16, -121, -128, 56, 99, 2, -4, 18, 58, 100, -32, 49, 110, -65, 98, 79, -51, -98, -69, 72, -101, -72, -8, 47, 40, -108, -92, -12, -113, -12, 101, -1, -4, 101, -72, -33, -24, 52, 113, -94, 25, -47, 83, 7, 16, 53, -42, 93, 84, 18, 37, 111, 74, -98, 30, -14, -78, 67, 102, -63, -73, 76, 65, 51, 49, 121, -109, -103, 45, -124, -69, -58, -42, -114, 77, 102, 68, -92, 68, 24, 54, -23, 7, 0, 7, -91, 114, 57, 104, 89, 123, -96, 37, 60, 83, -42, 53, 102, -16, -30, 107, 43, 41, -63, 58, -10, -89, -2, 26, 107, -106, -48, -43, 29, 80, 92, 66, 67, 22, 43, 28, 17, 75, -63, -51, 30, 23, -126, 5, -121, -28, -16, 51, -115, 49, -19, 4, 88, 107, -98, 68, -127, -17, -103, 30, -65, 117, -32, -126, 11, -117, 30, -100, 86, 95, -23, -11, -9, -21, 122, -2, 80, -22, -79, 93, -101, 30, -31, 115, 9, 0, 55, 10, 111, 80, -88, -82, 70, 9, -79, -47, 20, 79, -18, -21, 47, 87, 96, -90, -61, 90, 36, -109, -60, 86, 112, -33, -12, -46, -46, 126, 82, -118, 8, 65, 90, 49, 111, 32, -70, -96, 114, 78, 112, -32, -71, 31, -73, -103, 69, -6, 115, -23, 13, -73, -65, -2, 22, 52, 80, 105, 50, 34, 115, -70, -29, 77, 107, -46, -18, -91, -13, -32, 116, -29, 64, -83, -126, 119, -57, 71, -14, -70, -80, 127, -14, -16, -3, -120, -92, -51, 113, 86, 111, 100, -112, -46, 50, 124, 37, -96, -95, -104, 0, -107, -5, -64, -61, -3, -73, 10, -60, 41, 68, -12, 41, -74, 100, -90, -65, -120, -12, -80, 94, -29, -107, 111, 54, 71, 107, -37, 103, -116, -13, -25, -94, 110, 39, -27, -21, 94, 111, 47, 8, 51, -93, -79, 106, -120, -41, -87, -112, 75, -39, 111, -81, -18, 94, 101, -75, 73, -64, -100, 85, 51, 3, 119, 33, -86, -36, -116, -119, -53, 59, 17, 127, 94, 66, 105, 102, -103, -110, 119, 101, -21, 102, -108, 90, 68, 121, -113, 13, -71, -84, -30, 108, 47, -38, 13, 90, 54, 25, 99, -126, -44, -12, -127, -78, -74, 106, -103, -49, 124, -112, -76, -25, 118, -56, -63, 58, -63, -47, -57, -6, -3, 41, -26, -84, -125, 115, -122, 58, 12, 105, 60, 96, -35, 61, -109, 19, 39, -84, 99, 35, -68, -105, -118, -78, -32, -52, 108, 33, 29, -77, -100, -102, 92, 2, -58, 96, -10, -51, 26, -126, -74, -42, 99, 20, -109, 118, -89, 58, -94, -118, -35, -34, -94, -25, 16, 2, 51, -4, -93, -48, 47, -65, -22, 11, 66, 49, -21, -72, 126, -123, -70, -76, -37, -99, 72, -18, -109, 112, -88, -75, 122, 5, 19, -100, 109, -93, 30, 32, 31, 66, 113, -50, -127, -37, 90, 67, -116, -59, 123, -118, -53, -74, -65, 38, -45, -121, -107, -25, 119, -67, 28, 114, 67, -80, -114, 48, -45, 45, -48, 115, -17, -63, -63, -16, 29, -101, -76, 41, -31, -81, 52, 44, -27, 115, -46, 57, 122, -25, -96, 114, 37, 60, 100, -24, 108, 114, -104, -64, 31, -24, -77, -114, 42, -12, -1, -57, 16, 51, 112, 113, 98, 36, 29, -56, 23, 111, -127, 18, -41, -95, 4, 124, 93, -24, -28, 74, -38, -4, -118, 122, 100, -67, -120, 14, 49, 7, 85, -63, -70, 70, -78, -99, -22, 79, -27, -126, 63, -26, 20, -106, 7, -104, -110, -28, 0, -10, -82, 90, 114, -72, 84, 86, -11, 93, -27, -89, -28, -70, -24, 31, -128, 27, 60, -21, -22, -95, -19, -87, 7, -127, -65, -114, -103, -47, -14, 25, 71, 33, -13, 57, 89, -56, 16, -49, -91, 117, -10, 9, -81, 94, -88, -80, -7, 100, 27, 100, -123, -120, -115, 12, -119, -51, 26, -94, 30, -115, 59, -26, 46, -82, -97, 7, -10, 47, 86, 27, 36, -52, -91, 84, -85, -51, -124, 36, -78, 31, 8, -73, 39, 22, 68, 48, 99, -34, 82, 1, -21, 13, 103, -103, 59, -121, 33, -78, 54, -9, 77, -37, 68, 114, -81, 111, -64, -77, 19, -14, 82, -100, 41, -7, 50, -19, -87, 21, 76, 123, -106, -73, 8, 126, -47, -61, -123, 114, -11, 59, -23, -61, -106, -83, -75, -59, -100, -11, -8, 48, 103, -54, 76, 17, 67, -2, 126, 108, -109, 74, 103, -87, -126, -17, -89, -45, 51, -84, -59, -88, 104, 46, -21, 126, 92, 33, -60, 120, -106, 60, 40, 126, -121, -12, 15, 74, 114, 13, 55, -123, -40, 30, -81, -38, -114, -42, 45, 65, 3, 114, 105, -21, 32, -43, -23, -4, 118, 45, -11, -116, -22, -99, -118, -15, 18, 25, -69, 4, -89, 114, 10, -1, 17, 57, 89, 31, -113, 6, -32, 18, -8, -55, 125, -104, 30, -25, 21, 20, -108, -118, 33, -2, -89, 43, 111, 57, -59, -85, -66, -20, -99, 72, 107, 46, 1, 68, -51, 16, -54, 45, -93, 66, 119, -96, 90, 21, 7, -17, -86, 28, -7, 75, -102, 33, -10, -118, -38, 59, -75, 24, -89, -46, -32, -110, -127, 97, 86, -50, -14, -96, 124, 21, 98, 115, 53, 61, 8, -67, -84, 50, 89, 38, -3, 115, -57, 116, 125, 33, 47, -78, -70, 87, 5, 26, 105, 6, -4, 64, 84, 110, 96, 80, 3, 67, 67, -72, 0, -52, -11, 44, 126, -50, -46, -4, -62, 25, -16, -65, -69, -97, -14, -11, 118, 119, -113, 96, -3, 11, 32, -47, -7, 0, -94, 124, -61, 101, -75, 67, -79, 42, -16, -80, 121, 66, 44, -69, -36, -100, -6, 23, -69, 108, -116, -78, 99, -101, -110, -32, 39, 50, 50, -96, -78, 84, -99, -10, 57, -46, -71, 107, 124, 41, -101, 117, -20, 71, -80, 72, 99, 43, -33, -98, 23, -21, -48, -5, 6, -30, 91, -83, -108, 13, -50, -57, -31, -21, 61, -101, 61, 118, -122, 57, 32, -95, 47, -116, 104, 95, 84, 75, 10, -77, 105, -94, 30, -70, 29, -92, 28, -8, -46, 49, -122, 32, 120, -25, -117, 53, 2, 72, 43, 8, 1, -53, 41, -80, -41, 17, -112, -85, -36, 26, -34, -58, 60, 124, 0, -39, -95, -100, 82, -13, 77, 88, -109, 69, -65, -98, -6, 66, 102, -90, -54, -25, -15, 116, 24, 73, 5, 40, 116, 98, -62, -45, -88, 127, -49, 40, -40, -16, 68, -86, 99, 18, -126, 118, -41, -62, -108, 82, -124, 122, 120, -50, -30, -23, -62, 122, -78, 72, 34, -89, 42, 100, -6, 82, 99, 73, -6, -68, -70, -66, -26, -99, 80, -23, -108, -88, 43, -88, 122, 47, -93, 114, 125, 5, -37, -64, -1, 14, -120, -95, 53, 50, -123, -81, 4, 105, 120, 126, -91, -78, -68, 11, -48, -115, 116, -28, -75, 31, 12, -81, -50, 47, -95, -52, -76, -4, 12, 51, -118, 20, 84, 63, -58, 90, 110, 74, 67, 103, 72, 104, -103, -124, -13, -23, -111, -24, 77, -58, -121, -38, -11, -42, -119, 22, 34, -66, -109, -82, 113, -99, 66, 70, 93, -120, 32, 75, 82, -29, 50, 26, -53, 76, 30, 62, -75, 48, -90, -125, 118, -82, -35, -20, 4, -26, -126, -90, 36, -107, -44, 22, -77, -106, -36, -112, -98, 124, 91, 112, -33, 14, 10, 42, -38, -88, -24, 15, 88, 15, 18, 79, 61, 111, -69, -63, -42, -67, -25, 122, -45, 59, 16, 6, 81, 108, 22, 111, 104, -15, 95, -57, 127, -23, 113, -39, 17, -38, 105, -22, 105, -5, -71, 38, -21, -12, 103, 65, 49, -50, 59, -124, -119, -52, 10, 90, -72, -96, 73, -95, 18, 40, -24, 17, -111, -38, 107, 34, 52, 84, -116, 29, -49, -59, -61, 58, 57, -86, -5, -21, -8, -73, -17, 1, 3, 122, -37, 59, -102, -92, 92, 44, 76, -59, -66, 93, 31, -87, -1, -45, 125, 12, 112, -52, 81, -77, -121, 11, -35, 2, 118, 85, 57, -27, -42, -68, -33, 49, 120, -6, 85, 84, -90, 33, -103, -28, -2, 56, 13, 125, -117, 10, 9, 123, 87, -37, -82, 94, 102, 11, -32, 92, -32, -102, -63, 54, -42, 33, -25, -50, -101, -68, -93, -63, 93, -68, 38, -37, 117, -77, -39, -128, 62, 98, 124, 21, -67, -86, -13, -93, 54, 83, 127, -106, 109, -63, 77, -60, 98, -76, 18, 125, -15, 53, -66, -50, 114, 100, 42, 103, -104, -125, 103, 86, 101, 99, -21, -93, -114, 94, -58, 68, 49, -58, 90, 31, 7, 39, 99, -23, 92, -11, -26, -51, -85, 36, 27, -99, 9, -59, -124, 33, -56, 107, -9, -82, 79, 98, -47, 93, 64, 23, 33, -15, 93, -5, -112, -28, -93, 115, 77, 127, -23, -77, -52, 20, 88, 103, 49, -31, -83, 53, -126, -11, 32, -7, 35, -17, -37, 116, -52, -101, 12, 109, 12, -23, -23, 29, 78, 12, 16, 27, 11, 121, 79, 87, 13, 39, 62, -66, -120, 107, 115, -118, -31, 20, 3, -124, -125, 94, 121, -48, 121, 5, -67, 5, 110, 38, -94, 60, -78, 51, -40, 61, 44, -89, 20, -70, 78, -45, -8, 86, -66, -20, 96, 31, -128, -29, 36, -125, -63, 29, -45, -70, -94, 17, 63, -112, -73, 98, 77, -22, 21, -91, -89, -63, -52, 60, -5, -102, -113, 116, 112, -51, -32, 80, 109, -32, -77, 17, -29, -12, -82, 55, 46, -48, -56, -19, -32, -1, -49, -83, 105, 100, -46, -111, -90, 30, 77, 33, 56, 92, 21, 40, -87, 117, -8, -106, -43, 43, 39, 57, -97, 85, -16, 77, -91, 56, -69, 6, -73, 10, 51, -95, -17, -122, -78, 21, 36, 127, -74, -35, 91, 76, -123, -124, 65, -2, -101, -105, -87, 66, 80, -55, 24, -64, -106, 61, 120, -47, -61, -81, 92, 119, -48, -53, 125, 2, 96, 33, 1, -106, 126, -36, 98, -124, -31, 36, 2, -4, 59, 43, -66, 11, 116, 86, 75, -117, 20, 67, -36, 87, 114, -72, 78, -61, 3, 75, 69, -29, -19, -57, -6, -21, 35, -36, -17, -124, -128, 113, 0, 59, 29, 63, -58, 17, 21, -111, 28, -87, 84, 121, -127, 71, -79, 79, -118, 53, 27, 79, -104, -120, -106, 18, -13, 58, 111, 99, 62, 111, 84, -65, 43, -15, 126, 113, -125, 19, -125, 31, 61, 87, 24, 62, 30, 74, 13, 40, -1, -88, -8, 23, -80, 14, -86, 36, -56, -103, 7, -121, -120, -37, -58, 51, 77, -60, 37, 80, 87, 40, -17, 20, -1, -120, -46, -98, 82, 96, 70, -47, -120, -66, 104, -71, 77, -110, 93, -107, -85, -28, -100, -76, 63, -30, 103, 12, 38, 12, -36, -2, -76, 76, -110, 52, 84, -27, 82, 38, -59, 24, 119, -51, 87, 95, 6, 36, 114, -29, 57, -99, 71, 86, -47, 7, -72, -71, -109, 95, 69, -16, -35, 122, -68, -17, 46, -112, 84, 0, 54, -103, -104, 45, -25, 111, 12, 109, 19, -2, -47, -51, 28, -104, -93, 109, 31, -37, -90, 51, -70, 108, -93, 23, 102, -33, -121, 20, -17, 91, -108, -91, 117, -84, 82, -36, -100, -34, -55, 47, 93, 26, 124, -7, 51, -97, -26, -46, -5, 13, -123, 53, -7, -88, -51, -33, 7, -44, 115, 118, -81, -121, -101, -92, -77, 109, 0, -49, -52, 74, 127, -87, -28, 123, 34, -105, -101, -120, -22, 22, 21, -17, -53, -114, 24, 24, -19, -97, 108, -32, -106, -100, -25, -79, -64, 27, -97, 65, 106, -21, 11, 105, 20, 111, 101, -74, -121, -128, -66, -15, 22, 84, 96, 97, 98, -8, -6, -48, 24, -26, 48, 46, 2, -104, 95, 67, 51, 126, 4, 29, -23, -113, 7, 125, 126, -20, -77, -123, -20, -14, -10, -126, -58, -41, 99, -88, 79, -35, -8, -25, 68, -87, -107, -58, -63, 117, -119, 116, 115, 13, 17, -35, 28, -104, -38, 27, 4, 14, 32, 112, -128, -105, 114, -58, -18, 86, -18, -67, -77, 103, 37, 119, -112, 58, -66, -47, 47, -57, -59, 35, 85, 86, -128, -15, 111, -38, -116, -13, 104, 45, -28, 104, 68, -42, -82, -78, -84, 29, -17, -32, 4, -108, -41, 20, 79, 21, 101, -2, 93, -86, -95, 50, -128, -95, -93, 111, -4, -80, -29, -28, 93, 71, -51, 33, -99, -5, 83, -54, -104, -62, 42, 28, -41, -127, -80, -90, 23, -107, 36, -12, -65, 70, -90, -64, 103, -55, -81, -29, -7, 18, 72, -42, -39, -107, 119, -9, 16, 74, 65, 41, -115, -21, -59, -28, -20, -10, 10, -125, 11, -82, -9, 75, 116, 29, -117, 92, 103, -70, -65, -32, 77, -121, 55, -90, -100, 46, 29, 45, -7, -34, -42, 6, 73, 27, 106, -74, -111, -12, -71, 29, 34, 49, -24, 23, -50, -13, -13, -75, 45, 50, 22, -6, 58, -51, 33, 86, 123, -66, 3, -12, 29, 89, 122, -26, -11, 100, 28, 6, -40, 86, -93, 123, 7, 11, 18, 85, 126, -123, -117, 44, 55, 33, -90, -15, 110, 71, -56, 105, -122, 75, -34, 35, 37, -40, -119, -102, -67, 38, 32, 21, -4, 68, 16, -125, -49, -94, 88, -50, -89, 99, 122, 95, 4, -96, -48, -14, 104, 24, -36, 110, -28, 58, 17, -119, -110, 26, -93, -49, -64, 67, 101, 60, 7, -11, 63, 87, 24, 24, -91, 63, -5, -97, 30, -128, -65, 111, -14, -89, 7, 78, -107, 107, 8, 38, 116, 27, -63, -105, 106, 1, 91, 79, -66, -30, -59, 125, -71, 93, 21, -34, 28, -111, -3, -69, -111, 61, -86, 3, 100, 49, -46, 122, 29, 90, 32, 17, -11, 97, 41, -32, -29, 4, -81, 33, 102, -12, 30, -96, -47, -76, -2, 110, -59, 124, -87, -42, 57, -45, 89, 29, -124, -85, 23, 33, -122, -72, -77, -5, -103, 92, 91, -4, -32, -117, -99, -58, -1, 60, -26, 81, 112, 101, 63, -75, 97, 104, 11, 26, -69, -28, -73, -65, 16, 79, 97, 22, -121, -108, -111, -96, 112, 109, 29, -48, 120, 58, 22, -9, -10, 125, -56, -26, 98, -121, 27, 67, 111, -90, -35, -86, 11, 20, -22, -101, -29, -53, 49, -22, -33, 66, 11, -49, 47, -88, 31, 39, 98, -75, -97, -39, -78, -25, 63, -108, -17, -37, 87, -34, 1, -76, 9, -116, 73, 115, -89, -84, -66, 88, 23, 29, 27, -94, 108, -54, -54, 11, 114, -84, 64, -111, 5, 115, -8, -59, -121, 103, 32, 95, -58, -95, -109, 79, -82, 92, 66, -43, -119, -128, -82, 32, 29, 73, 66, 9, -109, -116, -108, -123, -72, 84, -106, 62, 71, 15, -125, 79, -10, 35, 46, 60, 68, 65, 11, 114, 30, -51, -56, 39, -51, -10, -57, 106, -65, -119, -13, -46, -107, 7, -40, -51, -36, -18, -117, -93, 125, -114, 114, -12, 49, 32, -80, -10, -30, 60, -24, -128, -119, 48, 39, -41, -90, 110, -63, -27, 119, 53, 56, -116, -68, -112, -39, 24, -2, -27, 60, -4, -13, 46, 112, -91, -49, -96, 27, 49, 92, -125, 49, 102, 52, -40, -67, 90, -58, -2, -64, -67, -77, 120, -55, -16, -120, 34, -120, 6, -121, 68, -126, -5, -13, 114, 32, 66, -109, -69, -13, 111, -66, -92, 85, 114, -4, -110, 77, 66, 17, -115, 127, 68, -123, -56, -76, -115, 106, -67, 19, 114, -127, 22, -19, -12, 8, -115, -74, 27, -56, 41, 11, 6, 77, -32, -7, -55, -13, -58, -117, -124, -45, -118, 72, -40, -46, 125, -27, -67, -70, 120, -81, -69, 14, 28, 48, -105, 41, 102, 50, 113, 16, -67, -9, -35, 30, 112, 39, -111, -74, 50, -107, 9, 61, 93, 97, -113, 90, -58, -52, -108, -65, -5, -48, 77, -105, -128, 100, 64, 102, 23, 49, -10, 84, -87, 84, -14, -103, -5, 3, -48, -83, 24, 89, 106, -10, 59, 122, -48, -127, -58, -27, -64, 66, 53, -114, 89, 53, 114, 26, 27, 9, -53, -110, -34, -12, 102, 80, 14, -31, -44, 94, 14, 108, 55, -7, -30, -14, -13, 51, -12, 57, -104, 52, -5, 77, 66, -43, 2, 53, 111, -99, -66, -70, -81, 28, 47, -107, -19, -67, -10, 65, -101, -123, 45, 82, -2, -112, -59, 113, 67, 57, 42, 91, -19, -90, 40, -80, -5, -86, 101, -22, -57, -93, 36, -9, 64, -45, 12, -83, 16, -125, 110, 43, -120, 27, -2, 6, 43, 67, -9, -18, -4, -95, -55, 105, -57, 113, -103, 66, -101, 126, -84, -29, -94, 81, 90, 98, -92, -26, -113, 53, -23, 125, -32, -15, 24, 94, 119, -60, 33, -18, 50, -99, 16, 124, -121, 87, 109, -96, 26, -119, -97, 70, -20, -63, 23, -58, -93, 60, 44, -78, -15, -106, -81, 81, 7, 71, 48, -1, -117, -47, 109, 62, -17, -3, 58, -10, -43, 39, 22, 111, 48, 53, 53, -100, 118, -51, -30, -103, -119, -113, -53, -6, -91, -6, -53, 44, -62, 123, -85, -51, -51, -103, -117, 60, 22, 69, -78, 107, -19, 72, 90, -99, -2, 16, -70, -12, 93, 28, 14, 102, 43, 89, -32, 80, -44, 43, -3, 22, 39, 40, 99, 116, 65, 111, 48, -40, 52, 98, -61, -95, 42, -98, -65, -88, 46, -7, 29, 11, -107, -85, -15, 65, -124, 81, 17, -40, -4, -114, 110, -93, 55, 82, -105, -8, 65, 71, 80, -11, 41, -108, 23, -44, -78, 86, -4, 96, -49, -103, -21, -28, -60, 92, -91, -55, 45, 55, 33, -87, 69, 16, -51, -4, -30, -28, 117, -93, -84, 69, 24, 85, 89, -81, -87, -117, -123, 38, 107, -44, 63, -42, 57, -124, -78, 94, -51, 95, 21, 110, -119, -37, -2, -42, 87, 96, 58, 76, -125, 102, 18, 28, 60, -21, 75, 101, -9, 81, 11, -30, -91, -53, 57, 94, -49, 107, 61, 28, 75, -46, 10, 84, 45, -119, -86, 5, 105, 100, -47, 109, 75, 99, 9, 7, -49, -44, -20, 70, -91, 120, -88, -53, -61, 97, -87, 18, 77, 102, -82, 24, -71, 56, -20, 102, 65, 22, -21, 43, -6, 61, 24, -59, 32, -95, 76, 111, -11, -71, 53, 27, -79, 94, 102, -12, 63, -113, -122, 12, 118, -76, -92, -81, 108, 16, -107, 46, -90, 1, -39, 33, -66, 113, 102, 94, -110, 51, 78, 7, 108, 3, -94, -99, -31, -120, 17, -95, -104, 23, 45, -114, 75, 82, -67, 55, -30, -46, -27, 9, 83, 62, -86, -111, 47, -112, 112, 65, 67, 62, -55, 47, -63, -21, 76, 35, -12, -35, 68, 12, 116, -15, 26, 63, -61, 87, -9, 38, -87, 92, -81, 125, 27, -39, -114, -54, -23, 126, -116, -83, 60, -43, 92, 126, 64, 41, 33, -76, -122, -27, 64, 123, 86, -38, 58, -102, -79, -79, 64, -37, -114, 111, -40, 41, -56, -26, 115, 49, -27, 127, 94, -95, -44, 59, -97, -107, -28, 64, -55, -22, -91, -118, -27, 124, -28, -96, -106, 22, -47, 86, 113, -33, 69, -55, -120, -115, 47, 124, 62, -108, 123, 29, -74, -48, -40, -43, -27, 60, -106, 46, -90, -69, 56, 12, -73, -99, 44, -51, 51, 125, -93, 36, -35, 104, 109, -27, 117, 28, -31, 52, 49, -35, -47, 103, 45, 41, -68, -110, -27, -46, 64, 11, 14, -7, -105, 69, 22, 67, -109, -55, 65, -74, 109, -98, -97, 90, 3, -108, -10, 101, 72, -89, -62, -103, -114, 111, 66, -53, -127, -89, 29, 65, 51, -85, -70, 74, 113, 80, 14, -124, -103, -49, -70, -122, -19, -39, 96, 112, -18, -41, 85, -74, -2, -105, -48, 13, -122, -110, 88, -121, -70, -11, 73, 109, 33, -125, 55, 18, 84, -59, 22, 109, 20, 80, 116, -127, -86, 84, 114, 24, -85, 71, 78, 42, 95, -98, -73, 101, -79, -113, 109, -21, 4, 54, -40, -91, 57, -113, 55, 13, -43, -51, -5, 105, -98, -17, 107, -56, -61, 93, 96, -17, 36, 46, -103, 3, 77, -48, -23, 126, -33, -42, -23, 99, -116, 65, -119, 69, 80, 64, -45, -91, -114, 78, -113, -84, -67, 122, -12, 0, 87, -44, 111, -5, -126, -120, 127, 79, -40, -24, 77, 55, 62, -74, 27, 74, 119, 36, 15, 72, -28, 98, 109, -14, 48, 124, 30, 109, 118, -110, -18, 77, -26, -35, -55, -23, -26, -56, -72, 62, 48, -122, -10, -18, -68, -111, -72, -76, 53, 71, 124, -103, 42, 105, 12, -38, 102, -86, -56, 92, -67, 54, 42, 35, -109, 115, -116, -7, -69, -59, -72, 107, -53, 46, -39, 7, 63, 17, 59, -12, -40, 55, 13, -126, 33, -103, -35, 7, -60, 37, -29, 1, -37, -115, -92, -18, -128, -79, 104, -69, -10, -96, -90, 65, 78, -1, -56, 13, -112, -124, -127, -23, 59, 14, -21, -36, 40, 72, 99, 108, -19, -57, -19, 72, -44, 17, -73, -43, 66, -97, 16, -72, -65, 55, 121, -115, -74, -62, 26, -57, -58, 27, 48, -127, -87, -101, -34, 81, 100, -63, 61, -47, 8, -86, -102, 93, 60, -47, -78, -2, -16, 66, 55, 47, -7, 48, 60, 48, 114, -42, 119, -72, 113, 39, -70, -102, 66, 24, 108, 38, 89, 41, 120, -30, 84, -110, -65, 16, -29, -15, -114, 83, -77, 69, 2, 45, -10, -66, -35, -24, 20, -44, 33, 5, 123, 91, 31, 61, -13, 11, -28, -52, -75, -36, 46, -119, -18, 109, 25, 81, -34, 39, 36, 18, -19, -90, -65, 99, -28, 28, -53, 120, 112, 108, -3, 107, 71, -100, 40, -70, 40, -116, 7, 93, -24, -75, 102, 86, -93, -1, 39, 1, -90, -53, -109, 19, -15, -46, -10, 85, 110, 66, 77, 94, 46, -54, 73, -10, -25, -14, 48, -113, -2, -73, 108, 103, -19, 82, 61, 16, -47, -27, -111, -9, 48, -91, -117, -94, -9, 1, 119, -26, -61, 69, -60, 114, -113, -114, -24, -10, 0, -104, 5, 126, -48, -15, 101, 61, -61, 35, -51, 20, -120, -34, -116, 56, 3, -105, 90, 123, 24, 82, -31, 92, 23, 37, 78, 38, 51, -74, -99, -77, -50, 34, -78, 30, -108, -105, -37, -41, 58, 40, 108, 66, -121, 120, -5, 10, -113, -43, 5, 39, -89, 102, 3, 62, 12, -47, -27, -65, 7, 2, -13, 86, -92, 37, -12, -72, 60, 80, 16, -9, -8, -4, -71, -1, -12, 52, -118, 3, -118, 15, -86, -79, -10, 46, 112, -126, 127, -43, -63, 7, 87, 52, -35, 123, -39, 81, -76, -106, 33, 68, 13, -102, -64, 70, 25, 52, -5, 35, -73, 5, -77, -31, 54, 41, -113, 38, 43, -113, 123, 108, 22, 82, 33, 115, 78, 122, 68, -126, -112, -26, 70, 29, 0, -122, -28, -103, 58, 95, 61, 113, -28, 112, -46, -102, 25, -30, 65, -60, -15, 60, -80, -121, 15, 81, 122, -35, 76, 62, -33, 92, -92, -91, -6, 36, -85, 94, 62, 101, 61, -5, 86, -95, -21, -88, -69, -124, 10, 124, -56, 123, 57, -8, -126, -56, -54, 124, 37, -106, 59, -124, 114, 95, -87, -20, 4, -44, -54, -62, -71, -121, 61, -113, -88, -88, -73, -28, -84, 66, -32, -12, 61, -103, 108, 64, -31, -74, 60, -122, -52, -9, -118, -65, -41, -77, 43, 91, 7, 118, -99, 64, 125, 90, 79, -90, -126, -121, 10, -82, 73, 106, 34, 6, -124, 14, -58, -27, 69, -125, -20, -111, -6, -10, -48, 81, 42, 124, 44, -79, 114, 73, 114, 111, 35, 65, -107, 37, 72, 31, 83, 17, 10, -11, -104, 14, -124, -34, 115, 73, -31, -33, 90, 92, 86, -85, 45, 0, -89, -38, 49, -103, -93, 35, -120, 71, -27, -98, -20, -83, 61, -64, 63, -57, 53, 87, 85, 57, -75, 73, 2, 23, -88, -35, -13, 126, 8, -96, -2, 47, -6, -80, 72, 30, 83, 80, -27, -72, 110, 81, -26, 44, -111, -91, 115, 71, 124, 73, 0, -79, 18, -125, 72, 58, -32, -69, 57, 104, -36, -73, 23, 86, -25, -33, -12, -69, -81, 89, -13, -98, 43, 89, 74, 60, 126, 61, 3, 122, 6, -124, -84, -104, -121, 116, 83, -25, -80, 12, -49, 12, 67, 102, -30, -85, -59, 87, -26, -12, 48, 89, 18, -37, 51, -36, -104, 49, -102, 27, 44, 32, 31, 88, 57, 38, 76, 12, -115, 124, -104, -36, 8, 91, -62, 107, -122, 7, 66, -20, 124, -14, -58, 14, 78, 121, 107, 102, 42, -123, 1, -42, 37, -95, -82, -34, 71, 123, 106, 85, 119, -126, -79, 0, 94, -12, -21, 100, 123, -83, -47, 119, 31, 23, 6, -19, 16, -15, -45, -70, -10, 85, 17, -101, 118, 63, -6, 61, 58, -28, 18, 50, -25, 68, -78, -59, -72, 29, -87, -77, 74, -6, -85, -23, -111, 49, 87, 33, -94, -86, 92, 24, 127, -19, 51, 117, -84, -83, 51, 103, 18, -59, 25, 121, -119, 75, -66, -63, -24, -25, -11, -78, 98, 32, 27, 115, -47, -14, 21, -13, 29, -15, -117, 28, 94, 62, 18, -118, 108, -59, 113, -2, 10, 10, -9, 20, -43, 53, 85, 61, -100, -54, 111, 126, 106, 11, 114, -69, 125, 7, 46, 26, 120, 57, -73, 86, -8, 73, 96, -28, -114, 82, 98, 24, -36, -39, -84, 50, -114, -126, -17, -86, -52, -33, -87, -73, 106, -101, -14, 103, 34, -95, 2, 26, 90, 57, -16, -46, 2, -48, 54, 16, -94, 24, -88, -1, 113, -43, -79, 127, -41, 32, -86, 35, 127, -45, 90, 105, -18, -51, 81, -112, -18, -45, 42, -56, -116, -102, 27, 14, -22, -47, -98, 13, 106, -58, -116, 91, 27, -67, 91, 114, 93, -123, 22, 93, -40, -16, 70, 70, 61, 23, 86, -85, 106, 0, -12, 118, 26, -113, 4, -124, -32, 34, 17, -54, 105, 29, -90, 4, 90, -127, -9, 56, -122, -115, 21, -34, -3, -37, -92, -69, 115, 122, -26, 93, -6, 90, 84, -108, 105, -40, -104, -54, 123, 42, 20, 100, -57, 58, -24, -94, 59, 95, 90, 65, 108, -17, -97, -22, 74, -61, 37, 61, -67, -117, 27, 55, 102, -17, 75, 79, 71, 100, -103, 66, 14, 46, 38, 85, -24, -113, 119, -92, 110, 81, 101, 91, -64, -123, -59, -117, -56, 106, 72, 6, 117, -29, -67, 91, 82, -119, 43, 26, 109, 68, -36, -5, -14, -125, -48, 91, -110, -56, 127, -128, -103, 100, 91, -38, 105, -96, -27, -78, -118, -83, 56, -128, 17, 117, 91, -29, 126, 6, 125, 107, -53, -38, -26, 61, -35, 55, 24, -17, 127, 23, -17, -104, -4, -53, -14, -27, -21, 87, 23, -10, -123, -49, -10, 22, -59, -47, 121, -61, 88, 119, -81, -93, -47, 21, 96, 46, -52, -7, -99, -53, -112, 12, -28, 12, 87, 86, 114, -61, 46, 9, 57, 51, 89, -81, -55, -98, 0, -62, -31, -40, -71, 16, -5, 10, -90, -36, -72, -14, 85, -43, 62, 101, 98, -94, -14, 57, 120, -28, 124, 38, 109, 53, -39, 70, 100, 34, 100, -27, 101, -58, 61, -98, 86, -71, 41, 124, 21, 97, -17, -22, -73, -83, -49, -103, -49, 65, 82, -57, -91, 79, 110, -109, 4, -57, 89, -23, 106, 62, 78, 79, -124, 11, 109, 90, 68, 22, 87, -39, -8, -58, 67, 47, -13, -109, 72, 66, 84, 26, -119, 122, -23, 119, -115, 110, -65, 102, -41, -87, 36, -91, 120, 40, 48, 101, 3, -11, -4, -38, 78, 116, 32, 18, 35, -109, 37, -21, 85, -7, -123, 94, -13, -17, 86, 0, -35, -107, -25, 52, -66, -117, 89, -74, 52, 9, -101, -73, 126, 23, 17, 77, 11, -79, -33, -82, -60, -124, 25, -103, -3, 31, 119, 113, -114, 77, -15, -21, 98, 88, -97, -96, 100, 120, -42, 24, 1, -14, 79, 0, -119, -32, -51, 21, 17, 44, 67, 85, 48, -35, 110, -83, 124, 101, -98, -118, 51, 16, -11, 21, -24, 20, 54, -52, 12, -116, 100, -115, -2, 51, 13, 8, -109, 90, -99, 36, 6, 96, -7, -74, -67, -25, -28, -71, -51, 2, -61, -128, -110, 56, 21, -5, -52, -53, 71, 88, -40, 44, 102, 86, -33, -13, -34, -13, -50, -5, -105, 84, -36, 17, -117, 25, 120, -17, 83, -59, 113, -106, -59, -124, 79, 91, -1, -101, -90, -58, 116, -2, 114, 90, -43, -46, -51, 51, 69, 27, -81, 92, -16, 11, -19, -5, -92, -26, 106, 119, 43, 91, -114, 113, 95, 93, 76, -34, 120, 114, 37, 108, -15, 23, 70, 70, 105, -108, -7, 46, 47, 40, 11, -97, -77, 120, 26, -40, -34, 4, -49, -118, -32, -35, 123, -65, -70, 71, 30, -77, 57, -61, -97, -86, 90, 102, 112, 68, 122, -22, -14, 41, -110, 125, 73, -58, 118, -29, 30, -44, 104, 109, -34, -56, -53, -39, 7, 5, -96, -91, 56, 90, -24, 88, -124, -61, 62, 117, -121, 56, -33, -7, -31, -15, -9, -86, 55, -19, 14, -43, 65, -10, -61, -96, 62, 14, -7, -59, -109, 26, -21, 76, -12, 83, 36, -8, -106, -30, -19, -99, -102, 76, 23, -5, -66, -114, 38, 117, -5, -76, -53, -68, 42, 14, -36, -24, -100, 86, 45, -81, -16, -104, 123, 100, 108, 31, -36, -126, -127, 74, -96, -101, 22, 55, 23, 84, 69, -67, 74, -64, -15, -107, -4, -101, 35, 89, 3, 63, 47, -80, 110, -97, -55, 106, -125, -75, 9, -33, -73, 11, -87, -41, 38, 64, -114, -67, 20, 83, -6, -34, -109, 107, -13, 16, -122, -106, -23, 9, 85, -104, 58, 68, -73, -125, 46, -70, -72, -73, 25, -17, 66, 67, 71, -23, 3, 85, 38, -105, 41, -95, -10, 60, -116, 105, -52, -109, -128, 53, 28, 85, 77, -42, 25, -124, -39, -57, -66, 17, -1, 88, -127, -63, 27, 72, 42, -98, 29, -47, -75, -58, -14, 43, -125, -2, 21, -49, 17, 21, -123, -82, -22, 82, 4, -124, 87, 94, -53, -107, -17, 74, 109, -16, -116, 8, -72, 54, 38, 86, -121, 92, -100, -7, 7, -97, 120, -100, -17, 9, 49, -12, 55, -100, -58, -68, -96, -99, -102, -21, -77, 9, -74, -96, 122, -62, 41, -78, 120, -49, -120, -128, -85, -91, -7, 51, -60, -15, 79, 51, 123, 1, -89, 50, 29, -18, 110, 61, 11, -120, -88, 62, 18, -34, 95, 12, 32, 8, 62, 25, 87, 71, 25, -125, 108, -110, 54, -80, 4, 5, 100, -1, -122, -117, -79, 35, -7, -96, -32, -123, -88, 9, 67, 58, 103, 34, -58, 8, -86, -123, -95, -126, 76, 58, -123, 56, 76, 59, 104, -48, -64, 76, 79, -57, 88, -127, 106, -47, -95, -53, -42, -55, 84, -102, -124, 59, 60, -54, -61, 103, -49, -28, 105, -101, -98, 110, 83, 107, 41, 60, -69, 105, 8, -117, -80, -32, -116, -101, 50, -83, -26, -120, -10, -70, -94, -6, 117, 95, 69, -71, 70, -108, 29, 47, -80, 60, 29, -125, 39, -58, 63, 98, -81, -56, 109, -32, 40, 121, -5, -38, -90, 97, -29, 29, -101, 5, -105, -112, -28, 92, -55, -86, 113, 103, 89, -95, 35, -10, -92, -54, 60, 100, -84, 108, -84, -102, -52, 84, -109, 71, -81, -70, 40, 18, 87, 67, -105, 110, 83, -4, 75, -99, 38, 60, -124, 0, 93, 39, 118, -127, 113, 51, 101, -99, 31, -111, -73, 107, 102, -53, 50, -107, 5, -38, 39, -36, -99, 62, -54, 112, -70, -107, -115, 97, 81, -111, -31, 46, 56, -41, 48, 41, -118, 21, 71, 41, 39, 126, 20, 13, -55, -58, 34, 78, 32, -55, -86, 61, -121, -11, 46, -62, 10, 59, -93, -36, 77, 4, -118, 5, 91, 58, -81, 102, -48, 118, 15, 119, 116, -92, 4, -66, -22, -90, -116, -117, -17, -73, 72, -10, 44, -10, 56, -74, -78, 91, 18, 127, -33, 29, 4, -69, -41, 51, -95, 39, 41, 48, 30, 30, 84, -94, 92, -65, -56, 104, -54, 55, -97, -110, -82, 75, 9, 102, -126, 59, 66, 20, 58, -95, -79, -66, -36, 9, 114, -3, -80, 27, -82, 79, -71, -126, 113, -107, -63, -70, 126, 11, 113, -99, 30, -97, 105, -89, -122, 107, 98, 72, -1, 28, 105, 49, 90, -58, -70, 76, 67, -22, -24, 113, -71, 33, 116, -85, 55, -75, -27, 53, 65, -42, 82, -33, -10, 59, 6, -4, 38, -24, -60, -90, -124, -83, 87, 94, -13, -111, 43, -73, -5, -109, -88, 53, 52, -100, 96, -21, -46, -59, -96, -109, 27, 115, -14, -111, 46, 120, 13, -43, -32, 81, -5, -28, 127, -46, -62, -14, -29, 109, 41, 94, -128, 82, 19, 53, 110, -13, -96, -64, 56, -63, -45, -44, -76, 69, -27, 98, 61, 115, -73, -99, 68, 50, 1, 67, -124, 68, -74, -25, 49, 95, -58, 50, 49, 89, -25, 32, -51, 7, 96, -123, 72, -76, -39, 124, 121, 63, 95, 55, 50, -106, 84, -10, 73, -42, -70, 77, -102, -16, -75, 75, -49, -5, -3, -127, -44, 100, 33, 33, -20, 1, 39, -76, 53, -128, -79, 47, 63, -112, -26, -15, -90, -70, 104, 111, 16, -94, 61, 42, 18, 114, -10, 97, -19, 115, 98, 65, 88, 3, -29, -60, -123, -118, -8, 58, -118, 41, -23, 74, 57, 79, -69, 96, -118, -93, 79, 26, -59, 12, -59, 87, -2, 59, 57, 107, 46, 27, 45, 6, -97, -112, 74, -92, -102, -61, 94, -92, 108, -56, 110, 38, -105, -86, 6, -95, -51, -43, 60, 19, 98, -127, -22, -32, 60, -93, -52, -22, 63, 121, 113, 94, -119, 59, -126, -93, 126, 96, -57, 107, -88, -74, 17, -64, -32, -105, -31, 45, -20, -99, -64, -50, -98, 43, 47, 90, 78, 123, -59, 13, 116, -74, -21, 125, 113, -19, -96, 112, -50, -25, 91, -10, 29, -20, 54, 125, 3, -104, 43, 111, -75, 107, -66, -44, 22, 109, -82, -27, 104, -13, 114, 92, 41, -34, 89, 27, 75, 121, 11, -103, -32, -26, 16, 126, 82, -58, 123, -43, -34, 38, -60, 20, 18, 2, 104, -88, -17, -106, 13, -41, 10, 0, -77, -77, 94, -116, 78, 41, -123, -39, 67, -26, 63, -45, -28, 17, 25, -33, 102, 120, -122, -85, 12, 24, 45, -12, 64, -99, 10, -50, -12, -108, 78, 40, -56, 44, 52, -106, -43, 58, -16, -104, -96, -81, -21, 4, 65, -123, 99, 39, 125, 105, 82, 9, 1, 0, 125, -62, 29, 7, 16, -111, 28, -34, 57, 100, -118, -18, 122, -33, -88, -22, -8, -56, 26, 99, 76, -37, 104, 47, -126, 101, 25, 85, -18, -102, -43, -21, -36, 114, 115, 108, -125, 15, -54, 61, -13, -44, -85, -19, 52, -45, 88, -84, 27, -14, -113, -25, 77, 120, -106, 79, 93, 47, 36, -52, 74, 121, 55, -90, 107, 42, -109, 111, -71, -35, 44, 44, 50, 87, -102, -26, -86, 114, 18, 69, -28, 33, -84, -79, 25, -62, -128, -9, 114, 37, 67, 60, 30, -6, 98, 10, -91, 117, -7, -34, -45, -91, -117, -123, 124, -91, -21, -90, -105, 125, 107, -5, 30, -105, 44, -72, -39, 44, 47, -53, -47, -14, -121, 112, 108, 106, -6, -111, 95, 115, -16, -78, -104, -5, -73, -108, 32, 34, -70, 55, 31, -91, -78, -66, -68, 94, -10, 21, 10, -91, 97, 92, 23, 104, 76, 3, 82, -58, 21, 50, -71, -123, 100, -47, 0, -100, -27, -96, 62, 31, 87, -34, 68, -119, 28, -128, 103, -110, 21, -15, -73, -10, -51, 78, -33, -103, -47, -79, -33, 102, 99, 24, 107, 72, 105, -21, 100, -50, 11, 34, 109, -30, -128, 49, -21, 28, 49, -46, 46, -57, 68, 101, 61, -111, 51, -100, -85, -123, -50, 10, 107, -79, -93, 87, 121, -116, -62, 93, -37, 78, 0, -56, -80, 0, 122, 28, -99, 43, 110, 75, 114, 50, 49, 48, 68, -28, 76, 111, -23, -102, -7, -43, -52, 28, -84, -59, 41, -18, -93, -124, -68, 35, -52, -19, -93, -58, -119, -64, 114, 119, -116, 100, 42, 61, 20, -18, -95, -31, -35, 11, -5, 86, 96, 71, -13, -116, -115, -100, -6, -80, -96, 55, 83, -20, -92, 118, 51, -83, -73, 37, -92, -61, 9, 78, -128, -98, -68, -95, -1, 25, 44, 122, -16, 12, 66, 99, 24, 79, 127, -109, 127, -97, 74, 82, 11, 110, 72, -66, -101, 127, 99, -65, -62, -19, -114, -62, 11, -54, -28, -118, 100, -112, -124, -44, 29, 70, -73, -75, 21, -74, -56, 20, -43, -110, -26, 96, -128, -81, -97, -101, -82, -126, -37, -15, -17, -23, 51, 122, 51, -105, -124, 23, -88, -119, 107, 69, 79, -94, 122, -27, -40, -61, 121, 45, -43, -32, 14, -42, 15, 45, -15, 61, 47, 76, -82, -97, -75, 98, -103, 105, 121, -98, 0, -95, -89, -20, 102, 118, 14, 97, -37, 103, -92, -43, 20, -7, 53, -94, 79, -60, 79, -63, -127, -1, -115, -80, 30, -61, -110, 55, -84, -117, 85, 44, -83, 124, -104, -109, 115, 39, 116, -50, 14, -104, 35, -94, 18, -40, -59, -31, 28, -108, 34, 30, 19, 48, 78, -79, 115, 96, 105, -97, 107, 62, 75, -104, 59, 100, -84, 46, 11, -96, 124, -103, -71, 32, -69, 75, 120, 0, -84, 21, 21, 79, -77, -88, -1, -127, -38, -14, 97, -61, 17, 76, -127, -36, 101, 60, -64, -111, -22, 75, -79, -25, 100, -22, -121, -96, -75, 127, 32, -30, 20, -75, -79, 71, -34, 48, 72, 56, -94, 41, 123, 51, -10, 124, -113, -37, 57, -48, -20, -93, -101, 29, 10, -128, -120, 17, -96, -67, 17, 64, 31, -91, 118, 80, 109, -44, 0, 53, -116, 34, -33, -121, -43, 85, -125, -27, -80, 60, 53, 28, 96, 80, -71, -22, 80, -63, 124, 112, -1, 13, 49, -98, 50, 39, 111, 31, 123, -17, -43, -121, -110, 52, -114, -25, 9, -111, 76, 57, 78, 1, -43, 46, -46, 14, -104, -94, 80, -108, -109, -49, 33, 68, -19, -44, -21, -36, 115, -26, 76, -56, -19, 94, 124, -5, -59, 5, 12, -110, -66, -38, 19, 19, -120, 101, -94, -95, -120, 114, -75, -101, -63, 87, 95, 46, -85, -54, -117, -98, 48, 87, -25, -99, 53, -29, 24, 122, 105, -92, -116, -89, -1, 32, 59, 7, 5, 93, 40, 13, 79, 94, 40, -112, 53, 7, 62, 96, 81, 73, 126, 1, 32, -27, 30, -43, 73, -74, -48, 50, -37, -36, 89, 90, 124, 20, -31, 2, -15, -118, -113, -64, 104, 56, -48, 29, -65, -113, -3, -111, 88, -5, 18, -7, 97, -79, 78, 42, -25, -98, -36, 66, -5, -75, 28, -9, 74, 126, 121, -69, -120, -119, -4, 112, 65, 76, 13, -128, 91, -118, -111, 52, 5, 36, -83, -26, 85, 123, -112, -68, -102, -20, 127, 21, 34, 27, -116, -20, 25, -122, 39, 33, -113, -93, 17, 80, 112, -98, 80, 75, -88, 98, -1, 46, 6, 44, -108, -37, 40, -91, 23, 66, 17, 22, -41, -77, -78, -29, 31, 75, -23, -57, -19, -8, -22, 126, -56, -38, -99, -103, -90, -59, 123, 37, 115, 1, -46, -120, 92, 122, -83, -13, 60, 62, -118, -109, 114, -68, -10, 17, -121, 96, 88, -12, -40, -61, -13, 33, 29, 16, 58, 67, 85, 53, -23, 73, -74, 59, 81, -110, 53, 126, 5, -15, 60, 15, 4, 46, 75, 122, -64, 83, 90, -104, -57, -77, -37, 58, 84, 121, -54, 14, 60, -96, -61, -91, 105, -7, 96, 58, 11, 21, 56, -112, -122, -12, 32, 10, -93, -21, 5, -29, -66, -33, -5, 6, 18, 87, -64, -26, 80, 11, 116, 12, 43, -73, 50, 20, 48, 18, -50, -69, -88, -122, -52, -82, -6, 108, 57, 29, -41, -66, -128, 22, 29, -4, -100, -80, -45, -36, 22, -93, 103, 11, 47, 18, 66, -31, -90, -13, 116, -12, 46, -100, -6, 122, -54, 117, 102, -125, 18, -66, -63, 19, 84, 95, -113, 112, -113, -30, -52, 37, 5, -76, -80, -76, 70, 115, 22, 109, -26, 10, -31, -108, 38, 92, -113, 112, 81, 117, 116, -29, -77, -75, 118, -121, -108, -123, 119, -93, -25, -60, 73, 108, -8, 121, -95, -66, 108, 55, -85, -46, -63, 13, -25, 103, -23, -10, 87, -70, -21, 75, 29, 31, -127, 20, 38, -107, 25, 30, -71, -127, 98, -126, 109, -38, 123, -114, 24, 104, 69, 68, -70, -122, -47, 33, 109, 58, -105, 69, 116, 3, 16, 17, -94, 17, -91, 72, 39, 63, -26, 96, 64, -56, 98, 45, 34, 93, 60, -69, 69, 1, 127, -128, 8, -48, 33, -11, -118, 57, -70, 126, -68, 75, 15, -34, -36, 53, -90, -125, -12, 13, 99, -76, 85, 69, 97, -8, 35, 29, 51, -24, -97, 50, -24, 39, -126, -118, -100, -116, 67, -41, -118, 127, -94, 25, -35, -2, -50, 3, 2, 66, -112, -27, 118, 102, -85, 88, -34, 78, -11, -111, -74, 20, 67, 31, -69, 69, 41, -40, 81, -20, 47, 91, -21, 81, -12, 72, -49, 67, -53, 81, 5, -36, -73, -4, -62, -30, -44, 32, -80, 73, 49, -26, -34, -12, -123, 25, -71, 46, 113, -118, -102, 32, 101, 5, -15, -39, -51, 65, -100, 25, 18, 34, 117, 73, -98, -73, -85, -14, 87, -37, -69, 8, 66, 25, 124, 71, -77, -75, -10, -92, -65, 16, 69, -92, -106, -74, -3, -29, 119, 26, 124, 10, -68, 113, -45, -38, -88, -1, 76, 127, 90, -121, 7, 28, 33, 3, -28, 84, 56, 90, 120, 119, -22, 61, -101, 0, 116, 25, 100, 107, -77, 96, -11, -17, 82, 73, 73, 122, -56, 21, 122, -94, 28, 1, 63, -67, -123, -93, -111, 61, 125, -118, 53, -25, 71, 80, 104, 59, -23, 76, 39, 28, 44, -100, -117, -2, 101, 84, -7, -83, -23, -13, -48, -122, 116, -113, -61, 121, -78, -43, 55, -81, -33, -20, 22, -90, -68, -2, 98, 38, -54, 9, -62, 119, 37, -50, -11, 11, -94, 110, 56, 12, -31, -120, 18, -42, -105, 85, -49, -55, -86, -122, -8, 9, -14, -113, 48, 47, 13, 18, -43, 88, -101, 23, 79, 64, 101, -60, -53, -120, -77, -124, 20, 20, -116, -90, 106, -92, 123, -70, -19, -90, -64, 102, 47, 51, 117, -33, -30, 2, 113, 55, -38, -116, -50, -87, 77, -76, -18, -104, -68, 33, -100, 80, -75, -87, 118, -96, -51, 113, -38, 58, -105, 26, 32, 71, -51, 21, -90, 47, -104, -104, -26, -14, -92, 53, 28, 113, 105, -118, -118, -91, 43, -90, 117, 96, -49, 107, -128, 28, 92, -38, -41, 116, 117, 119, 59, -62, 13, 97, 114, 37, 121, -40, -105, -98, -115, 51, -113, 118, 61, -103, -101, -24, -64, -112, -55, 15, 123, -55, -84, 88, 36, 3, 76, 25, -6, 7, 91, -121, -24, 77, 44, -30, -90, 68, 0, -77, -9, 15, -86, -75, 41, -59, 29, 105, -42, 102, -8, -47, -80, 36, -87, 84, -89, 117, -19, 34, -4, -56, 41, 101, -106, -42, -57, -68, -102, 71, -17, 17, -42, 25, 70, 127, 95, -28, 104, -75, -54, -31, 6, -6, -123, 48, -50, -83, 37, 59, 79, -94, -124, -8, -121, -102, 78, -50, -42, 104, -107, 69, -6, -21, -33, -64, -21, -66, 36, -45, -13, 111, 52, 121, -23, 58, 41, 56, 103, -49, -13, 54, -15, -9, -82, -8, 17, 125, 70, 103, 101, 91, 45, -33, -58, -116, 32, 49, -54, -60, -123, 61, -77, 57, 54, 29, -13, -32, -43, -38, 47, 72, -112, -96, -64, -65, 24, 81, -68, -34, 57, -95, -71, -26, 1, -1, -14, -95, -79, 60, -27, -74, -7, 25, 111, -81, -74, -29, 15, 11, 61, -66, -45, 78, -34, 19, -115, 118, -27, -55, -44, -98, -22, 13, 4, 107, -115, 118, -116, -66, 50, -14, -12, -85, -117, -29, -38, -63, 70, 106, 76, 4, -88, -97, -46, 7, 51, -33, -3, -104, 40, 82, -74, -110, -33, 58, 126, -20, 48, -118, 42, -30, -4, -98, 13, 7, 2, 103, 72, -56, 81, 20, 76, 122, 52, -98, 1, -25, -3, 126, -1, -91, 80, 53, -72, -80, -17, -74, 28, -97, -64, -57, 1, 61, -27, -114, -60, 103, 117, -115, -80, 71, 33, 124, 65, -43, -101, -62, 60, 24, -64, -69, 62, -111, 112, 118, -63, -33, -84, 93, -2, -20, -92, 127, -87, 10, -115, -18, -15, -125, -5, 33, 74, -100, 30, 11, -14, 57, 77, -82, -47, -115, -22, -113, -98, -38, -123, -33, 58, -79, -67, -72, 30, -31, -72, 71, 107, -59, -75, -35, -56, 48, 126, -110, 77, 28, 29, -65, -43, -22, -19, 39, -8, 87, 54, 22, -78, 60, 118, 108, 109, -77, -92, 11, 20, -36, -45, 0, 34, 8, 93, 106, -71, 91, 125, -122, -8, 26, -59, 77, -123, 50, -12, -3, 10, -85, -109, 60, 103, -119, 40, 84, -68, 76, -32, 81, -87, 51, -47, 75, -69, -82, 53, -12, -119, 50, -6, 1, -51, 63, -49, -46, -14, 67, 79, 124, 110, 98, 56, 85, 108, -32, 42, -88, -84, -118, 121, -43, 61, -54, -96, 120, -8, 86, -19, 2, 8, 103, -125, 85, 39, -46, -89, -103, -106, 118, -107, -124, 89, 77, 90, 69, -83, 4, 109, -39, 14, 103, 47, -53, -79, 79, -61, 42, 37, 48, -84, -82, 24, -81, -125, -65, 2, -85, -40, 24, -95, -19, 28, 122, -70, -10, 63, -25, 122, 45, 64, 8, 20, -17, 83, 69, -65, -105, -17, 100, 71, 27, -110, -33, 75, -106, 30, -51, -63, 118, 101, -30, -29, 1, -35, 29, 120, -100, -124, 114, 73, 69, -5, -35, -76, -50, -93, -13, -27, 18, -40, -83, -82, -22, 12, 121, 0, -85, -58, 65, -95, -85, -92, 5, 44, 1, -94, 36, 29, -89, 23, -25, 108, -110, 68, -96, -32, 103, 20, 70, -6, 108, 115, 40, -42, -1, 33, 87, 42, 103, 24, 76, -110, 60, -47, 62, -67, -13, -29, 91, 26, 122, -62, 6, -116, -122, 39, -20, 110, -69, -78, -24, -89, -91, -112, -3, 37, 49, -44, -49, 24, 109, -101, 42, 41, -20, -24, 103, 96, 75, 66, -6, 69, -124, -127, 81, -118, 40, -66, 120, 99, -16, -32, -118, 22, -16, 7, -69, -95, 92, 10, 57, 73, 38, -29, -14, -110, 76, -39, 114, 23, -101, -19, -35, -97, -18, -82, -86, -106, -20, -94, 121, 93, 3, -125, -13, 115, 10, 46, -107, -26, -72, 78, -81, 94, -78, 34, 113, 126, 123, 99, 21, -105, -48, 114, -74, 62, -95, -32, 84, 13, 3, 77, -22, -122, 80, 93, 121, -37, 11, -114, 65, 68, 93, 113, 34, -113, 19, 19, -115, 14, -9, 34, 37, 71, 21, 92, 6, 54, -68, -38, -61, 63, -88, 46, 69, 120, 11, 63, -45, -105, 77, -107, 91, 42, -122, -3, 57, 25, -111, 70, -89, 8, -23, 77, -49, 126, 41, 85, 52, 101, -80, 119, 37, -40, 37, -22, -48, -79, -87, 36, -56, 119, 57, -93, 33, 63, 32, -37, -40, 49, -95, -1, -71, 10, -52, 9, 8, 117, -34, -68, 91, 14, -76, 0, 102, 89, 106, -73, -118, -108, 91, -46, -117, 20, -11, 44, -45, -106, -121, 43, 71, -87, -86, -127, 51, -9, 10, -68, -20, 104, -8, -57, -9, 44, 71, -35, 6, 50, 20, 16, 70, -17, 99, 81, -125, -40, -3, -42, -18, 5, -127, -74, 46, -84, -73, -31, 35, 65, 29, -113, 41, -106, -41, -96, 66, -98, -2, -56, 80, -110, 89, 22, 2, 60, -25, 5, -108, 101, 92, 3, -22, 93, 57, -104, -119, 112, -7, 44, 49, -105, 60, -38, -83, -109, -5, 111, -79, 121, -72, -126, -117, -111, 24, 13, 77, -128, -109, 97, 101, 111, -28, -49, 76, -99, -25, 86, -115, 96, 2, 62, 119, -66, -103, -92, -47, 20, -108, 3, 13, -52, 5, 24, -35, -99, -90, -86, -99, -71, -117, -126, -88, -16, -47, 116, 13, 56, 74, 27, 25, -51, -39, 16, 11, -14, 53, 93, -122, 73, -32, 19, -107, 101, -84, -14, -126, -46, 28, -96, 11, 39, -94, 51, -105, -12, 39, 37, -84, -14, -64, 69, 63, 25, -42, -54, -116, -117, -89, -110, 84, 7, 38, 105, -20, 82, -37, -17, -92, 119, 15, 47, 30, 49, -30, 54, -91, -119, -37, -46, -5, 27, -105, -70, -76, -19, 5, -64, -8, 44, -45, -52, -76, 121, -75, 32, 75, 16, -113, 111, 7, 30, 30, -90, -48, -128, 92, -11, -119, -73, 71, 5, 82, 95, 63, -122, -52, -60, -57, 69, 113, 26, -111, -91, 19, -57, 69, -34, 87, 85, -51, -33, -13, 107, 5, 67, 107, -31, -71, 116, 24, -128, -7, -22, 95, -71, -16, -84, -3, 55, 113, -18, -47, -126, 19, 100, -55, -39, -62, -95, -82, 15, 0, 33, -6, -123, -27, -27, -26, 30, -38, 126, 30, 83, -24, -2, -116, 88, 42, 10, 16, 27, 120, 97, 29, 12, 70, 103, 101, -120, -120, -109, 24, 8, 52, -110, 13, -103, -8, 115, 55, 82, 113, -42, 37, -39, 84, 50, -79, -2, -68, 65, -103, -76, 35, 54, 64, -23, 29, 37, -15, 37, 56, -119, -83, -19, -100, 58, 6, 20, 45, -66, -26, 30, 20, -117, 119, -24, 61, -87, 102, 121, 106, 127, -82, 13, 53, 110, 118, -45, 20, -24, 120, -52, -15, -90, 57, 13, 96, -64, -95, 14, -2, 7, -84, -110, 19, -92, -6, -48, -51, -32, -54, -73, -33, -8, 69, -108, -26, 59, -25, 122, -93, -32, -57, 21, 6, -128, -94, -26, -64, -60, 116, 62, 75, -95, 80, -34, -59, -54, 47, 18, 42, 121, 73, -119, -15, 14, -98, 87, -54, 5, 82, -19, 101, -103, -126, -21, -103, -91, 82, -38, -23, 70, -104, -76, 103, 105, 19, -84, -77, -62, 62, 94, -69, 8, 103, 44, -106, -123, 3, -32, 11, -43, 78, -16, -18, 80, 92, 8, 117, 46, 98, -34, -12, 122, 19, -36, 99, -90, 8, -105, -24, -57, 117, 35, 79, 92, -49, 101, 98, 82, -58, -19, -88, -108, 93, 22, 100, 57, -98, 90, -25, -128, -72, 92, 123, 75, -72, 94, 113, 64, 117, -39, -121, 106, 124, 86, 71, -53, 60, 41, -98, -126, -106, -58, -106, 115, 92, 122, 45, 123, 84, -108, 123, -115, 112, 118, 88, -88, 85, 74, 105, 74, -93, 112, 53, -96, 71, -4, -21, 3, -91, 9, 5, -69, 79, 27, -82, 44, 21, 91, 39, -22, 112, 34, -9, 96, 25, -49, -119, -18, -103, 114, -72, -67, 98, 109, -35, 41, -23, 72, -84, 14, -46, 49, 73, -95, -52, 120, 77, 98, 83, -12, -52, 67, -105, 67, 36, 48, -110, 45, -98, -84, 31, -42, -23, 1, -60, 70, -85, 45, 14, -41, -68, 96, -119, -123, -126, -43, 125, 79, -73, 81, -60, 3, 20, -37, -58, -72, -117, -39, 101, -87, 5, 4, -1, 110, -122, 67, 52, -79, -15, -62, 8, 45, -93, 17, 50, -91, 103, 48, 116, -98, 1, -72, 34, -107, 19, 104, -50, 30, -63, -77, 71, 70, 56, -57, 52, 62, -118, -24, 111, -5, 43, -9, -88, 78, -119, 91, 115, 112, 11, 103, -114, -116, -96, 48, -95, 51, 25, -17, -46, 90, 35, -103, 33, -37, -32, -43, -103, -21, 62, -120, 102, -23, -1, -113, -73, 8, 106, -86, -8, -11, -111, 7, 1, -79, -73, 34, 101, 80, -110, -73, 43, 53, -48, -52, -112, 49, 33, -87, -100, -33, -79, -126, 72, 48, -111, 127, -71, 123, -87, 49, -16, -69, -72, 113, -20, -16, 20, -47, -64, 38, 8, 107, -37, 89, -73, -21, 10, 89, 20, 38, -72, 69, 40, -127, -11, 58, -128, 46, 53, -86, -32, -90, -27, 24, -105, 81, -120, 43, -93, -55, -47, 43, -76, 44, 4, -20, -105, -114, -59, 43, 52, -3, -16, -35, -2, 102, -105, -1, 20, 76, 41, 116, 114, -114, 13, -118, 95, 21, 53, -126, 94, -121, 46, -109, 51, -78, -1, 75, -63, 68, -10, 117, -63, 103, -46, 64, 77, -23, -65, -31, -74, 104, -42, -88, 118, 99, -78, 85, -8, 104, 88, -41, 111, 6, -22, 34, 56, 105, -19, 121, 45, 100, 111, 110, 75, -63, 46, 24, 43, 109, 121, 97, 85, -49, -119, 75, -78, -68, 33, 43, -92, -7, -126, -109, 127, -20, 53, 55, -43, -93, 49, -126, -121, 32, 112, 82, 97, 31, -22, 12, 12, -29, -19, -30, 51, -9, -83, 101, 51, 78, 16, 87, -57, 18, 106, -58, 126, 31, 126, -45, 66, 47, -43, 73, -49, -58, 27, -80, 101, -123, 61, -15, -23, -86, 83, -100, 33, -127, -127, -44, 79, 18, -85, -105, -92, -107, -35, -93, 53, -37, -10, -9, -118, 76, -63, -39, -110, 92, 10, 119, 98, -57, -24, -53, -15, -68, -25, -109, -67, -24, -25, -116, 122, 19, -93, -97, 40, 1, -62, -35, 92, 56, 85, 103, 4, -106, -64, 22, 114, 74, 13, 84, -111, 118, -97, 3, -78, 6, 22, -17, 111, 125, -5, 105, 16, 31, -120, -71, -96, -54, 22, 124, -125, -21, 99, 7, 1, -92, -98, -12, 110, 43, -56, -128, 33, -24, 3, 83, 110, -103, -62, 93, -106, 62, 71, 39, -35, 79, 96, -3, -102, -10, -7, -99, 98, -35, 36, -29, 1, 66, 87, -17, -18, -96, -17, -113, 8, 114, 99, -10, -117, -91, -44, -94, 99, -101, 73, -64, 106, 41, 61, -124, -97, -73, -95, -127, 20, 70, -27, -107, 8, -68, 4, 118, -36, 116, -122, 100, 102, 105, -37, 114, -114, 47, -108, 114, 74, 93, -78, 52, 6, 112, 57, 37, -89, 90, 39, 59, 32, -116, 80, -87, -56, -44, -97, 37, -56, -91, 9, -81, -114, 100, -95, -99, 19, -75, -113, -35, -110, -63, -110, 24, -79, 75, -67, -40, 37, 100, -109, -58, 112, 99, -17, -71, -72, 14, 94, 0, 52, -25, 47, 66, -52, 80, 95, 95, -123, 110, -67, -105, -80, -49, 47, -31, -102, 109, 58, 63, 81, 77, -123, 66, 49, -12, 123, 105, -125, 89, -23, 55, -64, -103, -7, 12, 105, -39, -20, 111, -57, 41, -122, -9, 120, 54, 89, -110, 35, 19, 81, -12, -32, 87, -74, -111, -53, -79, 122, -50, -118, -28, -123, -53, -3, -1, 87, -26, 88, -61, -43, -97, 108, -36, 23, 100, -110, -16, 118, 53, -125, 72, -87, -29, 31, -32, -11, 106, 17, -17, -71, 28, 83, -66, 103, -48, 61, 62, 55, 21, -126, -116, 53, 110, -24, -52, 83, -6, 60, 73, -81, 63, 17, -39, -94, -80, 57, 23, -101, -54, -121, -44, 102, 90, 18, 77, -85, -48, 12, 98, 101, 14, 110, 26, -4, -41, 102, -49, 81, 34, -103, -127, -31, 42, -38, 4, 91, -109, -101, 118, -35, -94, -54, -60, 125, 92, -111, -88, -84, 29, -118, -110, -85, 120, 44, 40, -49, 19, 119, -95, -75, -112, -94, 23, 59, -4, -101, 22, 15, -74, 12, 108, -39, 86, -80, -42, 50, -62, -2, 95, 95, 8, 113, -117, 0, 29, 51, 80, -80, 42, 113, -26, 59, -109, 125, -10, 15, -104, -116, -98, -50, 24, -118, 39, -18, -69, 125, -96, -3, -5, 127, -36, -125, 112, -25, 4, 14, -102, -44, 62, 69, -59, -92, 0, -40, -95, 118, 103, -71, -126, -123, 8, 26, -113, -81, -120, -54, -83, -88, 71, 40, -88, -92, 44, -104, 11, -80, 38, 38, 4, -27, -21, 73, 9, 107, -95, 43, 97, -120, 100, 99, -115, -20, -3, -100, 28, 5, -25, 73, 45, -82, -15, 85, -46, -99, 110, 94, -51, 20, 4, 81, 121, 111, 26, 3, 90, 59, -82, 59, 67, -110, 30, 80, -1, -101, 109, -101, 32, -44, 100, -51, 2, -43, -93, 85, -13, -111, 51, 64, 37, -73, 18, 31, -90, -84, -94, -128, 104, -48, 59, 43, -30, -39, -4, 97, -12, -23, 124, -108, 61, 96, -31, -65, -74, 4, -108, 41, 21, 71, -23, -69, 126, 123, 90, -92, -88, 124, -92, -112, -52, 95, 59, 46, -72, -73, 16, 44, 32, 12, 64, -35, -19, -94, 29, 35, 38, 49, -52, -68, -7, 53, -9, -9, 49, -47, 28, 89, -51, 64, 105, 25, 32, 36, -57, 88, 92, 87, 5, -4, -28, -59, 90, 81, -25, -9, -12, -114, -88, 64, -54, 33, -11, 65, -103, -90, -110, 53, 127, -33, -11, 104, 120, -107, 13, -65, 110, -23, -105, -13, 101, -5, 56, 63, -52, -96, -74, 64, -82, -33, 0, -8, -128, 117, -71, -103, -100, -53, 78, -101, 42, -60, -124, 34, -39, 17, 97, -57, 122, 120, 58, 95, -13, -13, 31, 63, 19, 85, -1, 65, -76, 127, -71, -75, 117, -14, -50, -111, 61, -99, -84, -25, -31, -80, -119, 58, 65, 106, -126, 59, 99, 60, 27, -42, -81, -70, -106, 66, -113, 21, 3, -60, 21, 60, -7, 10, -82, 71, 27, 107, 100, 71, -46, -59, 120, -37, -128, 57, -58, -126, -11, -87, 62, -112, -1, 110, -54, 21, 48, -39, -85, -76, 29, 64, 112, -106, -54, -97, 94, 101, -118, 66, 44, -35, -120, 36, 56, -120, -34, 126, -118, 83, -89, 72, 99, 39, 54, -83, -68, -25, 6, -25, 27, -92, -89, 11, -70, -15, 42, -104, -42, 53, 91, -125, -110, 99, 39, 74, 107, -123, 73, 117, 88, 112, 61, 59, 23, -12, 104, 84, 91, -17, -69, -10, 19, -29, -127, 77, 84, 44, 102, -85, -31, 65, -82, -13, 36, 85, -67, 15, 91, -122, 4, 51, 119, -63, -17, 14, 53, -41, -30, 16, 70, 30, -122, -39, -127, -120, -89, 85, 52, -115, -128, -107, 78, -82, 8, -14, -124, 69, -127, 95, 76, 5, 18, 67, 70, -127, -47, -4, -39, 52, -116, -97, -46, -109, -7, -45, -101, 32, -88, 79, 45, -87, 100, -5, -41, -20, 109, -37, -79, 110, -70, 125, -13, 77, 64, -71, 78, -110, 53, -89, 70, 66, -57, -104, 85, 64, -21, 112, -32, 19, 63, -115, 60, 35, 8, -108, -113, -11, -17, -64, -29, 42, -66, 86, -9, 126, -113, -59, -112, 69, -19, 86, 7, 52, 110, -36, -12, -39, -52, 84, 109, -117, 97, 41, 46, -23, 61, 61, 94, -83, 125, -63, 87, -69, -105, -50, -70, -90, 19, -54, 107, -128, -95, -14, 52, -113, 78, -88, -23, -102, 124, -42, -91, 93, 127, 83, -58, 61, 16, -92, 106, 14, -27, 65, 73, -4, -113, -125, 35, 34, -50, 14, 35, -17, -127, -41, -2, 79, 0, 103, 106, -4, -67, -113, -38, -67, 99, 32, 122, -13, 69, 100, -127, -86, 37, 75, 39, 52, 78, -54, -42, -100, 88, 121, 11, 89, -47, -118, 41, 81, 113, 19, -51, -81, 34, 39, -20, 5, -56, -26, 121, -115, -54, 122, -73, 111, 69, 94, 35, 20, -88, 121, 48, -127, 115, -68, 90, -60, -58, 3, -107, -73, -106, -30, -26, 57, -118, 82, -66, -46, -72, -73, -33, 2, -78, 22, -15, 119, -11, -108, 11, 29, -114, -68, 30, -127, -8, -7, -59, 62, 124, -38, 117, -109, 60, -36, 76, 70, -82, -118, -104, -25, -62, -9, 105, -12, -114, -37, -21, 3, -17, 119, -96, -3, -77, 63, -2, 43, -72, 67, -23, -76, -99, -34, -57, 90, 58, -109, 32, 105, -98, 57, -48, -32, -80, -71, 84, -66, 20, -65, 65, -124, -74, 98, 1, -23, 33, -128, -108, 89, 67, -3, -115, 97, 92, -43, 59, 22, -24, -37, -1, 6, -108, 79, 102, -59, -119, 58, 3, 29, 122, -59, 33, -80, -89, -93, 26, 72, -93, 46, 33, 102, -84, 46, 71, -120, -125, 2, 30, -20, 94, -98, 114, 114, 109, 89, -73, 118, 19, 59, 20, 13, -128, -75, 62, -89, -40, -40, 111, -5, -122, 16, -30, -78, -66, -87, -70, -62, 44, 89, 46, 10, 119, 32, -4, 100, -7, 52, 91, -115, -17, -17, 26, -17, 36, -40, 22, 125, 48, 5, -8, 55, -107, 90, 105, -45, -124, -92, 21, 48, 125, -61, -70, 116, 100, 54, 88, -35, -22, 51, -22, 89, -94, -123, -56, 71, -35, 94, 68, -114, -29, -68, 69, -8, -105, 46, 76, -101, 82, -31, 75, 79, 37, -123, 67, 9, 59, 28, 102, -90, -49, -47, 127, -14, -42, -56, -71, 51, -90, 125, 65, 10, -71, 6, -126, -48, -75, 78, -21, -121, -80, -74, 87, 85, -69, 26, -34, 119, -74, -60, -99, 6, 21, -100, 120, 107, -28, -79, 31, 11, -82, -32, -107, -25, 103, -105, 56, -100, 102, -93, -93, -106, -38, 122, 107, 21, 21, -55, 12, 75, 13, 41, -47, -93, 70, -55, -114, -86, -6, 45, 53, 40, -114, 74, -112, 117, 98, 72, -111, 72, 107, -76, 94, -59, -81, 73, 91, 68, -110, -25, 15, 31, -111, 97, 66, 87, -86, 81, -127, 37, -2, 55, -51, 12, 1, -35, 1, -29, -91, 18, -85, -111, 71, -119, -42, 118, 82, -79, 58, 100, 25, -55, 4, 42, -86, -58, 1, -43, -105, 2, 122, 22, -71, -57, -94, 59, 37, 36, -98, 74, -74, -54, 91, 125, -45, -78, 115, -90, -29, 45, -118, 124, 119, 14, 38, -95, 85, -89, -10, 108, 42, -16, 2, 99, 56, 37, 30, -35, -55, 61, -89, -1, -121, -125, -3, -38, -75, -16, 0, 24, -98, 11, 21, -107, -103, -69, -74, 110, -29, 45, 91, -115, -99, -35, 112, 85, -126, 15, -78, -53, -52, -38, 75, -45, -35, -56, 45, 18, 56, -82, -86, 86, 57, 63, 107, 82, 123, -94, 65, -34, 79, 28, -21, 108, 121, -37, 66, 124, 106, 116, -57, -74, -50, -110, 9, 43, -38, -73, -67, -109, -27, -24, 105, -98, -89, 85, 112, -94, 119, 49, 0, 70, -51, 107, 50, -57, -57, -12, -61, -79, -23, 10, -24, 55, 29, 113, -29, 119, -88, 32, -118, 13, -120, 116, 43, -80, 73, 28, -46, 64, -51, 83, 6, 27, 62, -72, 98, -123, 45, -91, -73, -106, 47, 31, 77, -52, 16, -80, -60, 57, 81, -50, -58, 89, -62, 114, -119, -117, 14, -36, 75, 91, -81, -47, -10, 109, 10, -40, 115, -73, -3, -86, -51, -83, 73, -102, -7, -39, -53, 61, -110, -100, -116, -39, 117, -50, -53, 127, -38, 89, -37, -91, 52, 10, -9, -85, -9, -127, 3, -22, -72, -127, 20, 5, -82, -35, 31, 39, 55, 106, -27, 73, -122, -15, -94, 124, 63, -19, 123, -103, -58, -42, -65, 123, 96, 54, -90, -41, 55, 41, 66, 111, 42, -42, -12, 88, 52, -109, 0, -21, 126, 101, -76, -124, -42, -41, -128, -107, 68, 123, -81, -117, -47, -18, -122, -79, -92, -84, 9, 91, 85, -53, 74, 0, 33, -66, -40, -43, -47, 88, 64, -49, 61, 117, -44, -109, -52, -44, -87, -112, -48, -40, -101, 33, 70, -95, 83, 106, -51, -36, 69, -93, 39, 15, 35, -56, 77, 123, 30, -98, 84, -34, -18, 17, -45, 66, 37, 31, -106, 78, 48, -26, -90, 75, -120, 108, 109, 91, 86, -70, -73, 27, -35, 94, -86, -128, -90, 119, 124, 68, -107, 80, -93, 3, -31, -10, -59, -122, -106, -36, 84, 70, 66, 122, 17, 74, 102, -2, 37, 60, 57, 92, -41, -106, 58, 1, -105, 97, -8, -109, 37, 14, 99, 72, -111, -60, -65, -41, -53, -43, 51, -97, -101, -11, -102, 44, -64, -128, -85, 101, 61, 100, 66, -108, 122, -4, 22, -111, -35, -114, -92, -125, 28, -121, 75, 46, -52, -118, -123, 23, -33, 56, 54, -6, -83, 80, -89, -19, 81, -46, -45, 14, -74, -107, 34, -80, 17, -72, -62, 111, -57, -26, 114, 99, -18, 61, 17, 58, 72, 22, -47, -89, -50, -121, 34, -4, 88, 73, 105, 41, -101, -68, -73, -47, -47, 89, 1, 99, -110, 67, 82, -39, -86, 68, -68, 24, 1, 78, -46, -55, -28, 35, -15, 51, 42, -109, -81, 2, 92, -104, -85, 119, -43, -30, -56, 38, -68, 73, 9, -50, 13, -37, 39, 55, -97, 99, -49, 33, 49, 33, 106, -106, -60, -37, 73, 110, -18, 120, -15, -54, -112, 28, -63, -27, 127, 9, -116, -69, -45, 21, 9, 96, 113, -80, 23, -112, -109, 102, 49, 69, 7, 28, 91, 75, 119, 36, 57, -26, 28, -86, 48, 44, 71, 114, -110, 70, -5, -98, -127, 78, 51, 10, 46, 36, 58, -59, 53, 77, -85, -26, 18, 50, -126, -19, -3, 122, -111, -73, -32, 45, -31, -112, -38, -88, -126, -20, 110, -2, 10, 111, -52, -67, -7, 123, 98, -77, -64, 23, -127, -20, 125, 19, -98, -128, -127, 28, 122, -110, 83, -38, 64, -76, -22, -102, -35, -19, 6, -53, 107, -112, -69, -73, -51, 52, -78, -81, 104, -13, 70, 105, 95, 68, -4, 125, 68, -3, 25, 62, 16, -20, -104, -48, 33, 2, -22, 126, 111, 112, -55, 90, -128, 4, -110, -51, -71, -60, -3, -95, 55, -61, -118, 22, -121, 6, 20, 75, -124, -83, 9, 20, 26, 33, 100, -69, -92, -50, -71, -109, -66, 2, 110, -66, -121, -128, 11, -64, -60, -120, -31, 124, -52, -21, 18, -45, 113, -90, -97, 117, -44, 40, 9, 110, -54, -19, -87, -18, 59, -30, 1, 121, 100, -17, -73, 107, -17, 67, -85, 52, 75, 12, 48, -105, 119, -62, -21, 105, -23, 10, 94, 61, -78, -24, 43, -4, 85, 84, 106, 17, -74, -20, 10, -102, 91, 66, -122, -53, 5, -79, 127, -48, 62, 47, -24, 53, 113, 83, 30, -38, -35, -3, -105, 15, 101, 66, -116, 58, 22, 118, -53, 76, -30, 86, 103, -66, 24, 109, 9, -99, -98, 8, -19, 92, -73, 85, 18, -88, 40, -80, 3, -123, 45, 26, 21, 18, -35, 33, -51, 115, 23, 24, 64, 122, -18, 39, -72, -122, 20, 65, -93, 50, -55, 17, 15, 0, -26, -95, 40, -113, -47, -85, -108, 127, 70, 41, 17, -93, -54, 94, -106, 98, -9, 86, 92, 101, -3, -108, 108, -111, 85, -113, 68, -98, 32, -45, 30, -121, -12, -58, -106, 69, -14, -86, 68, -72, 84, -42, -37, -98, -76, -15, -128, 43, -56, 92, 17, 69, 112, -3, 87, 69, 12, 27, 99, -83, 110, 1, -76, -30, 72, -54, -89, -70, -12, 108, -14, -56, -62, 77, -25, -10, -66, -25, -94, 6, -60, 51, -52, -76, -80, -93, 122, 60, 62, 93, 105, 44, -33, -99, -114, -89, -25, -75, -31, 92, -95, 83, -92, -29, 32, 11, 90, 94, 115, 124, -27, -73, 47, 49, -21, 95, 84, -27, 27, 18, -61, 5, -66, 34, 34, -52, 73, -118, 1, -86, 102, 35, 125, -118, -122, 29, 22, 96, -5, 9, 92, 96, 64, 11, 17, -85, -22, -27, 17, -122, 119, 84, 11, -75, -10, -83, 1, -65, -73, -125, -23, -99, 38, -26, -88, 44, -125, 62, 13, -2, -57, -23, -33, -121, 117, 112, -78, -33, -42, 67, -27, -51, 23, 112, 3, -115, -98, -124, -52, -43, -121, 53, -13, 45, -101, 27, -38, -98, -39, 103, 29, 32, -48, 124, 39, -59, 108, 89, 37, -62, 29, -118, 16, -76, 123, -109, -62, -103, -105, 14, -18, -97, -60, 97, 76, -33, -4, -90, -2, 85, -115, -101, -11, -34, -105, -100, 35, -125, 118, -56, -58, 19, -45, 86, 71, -50, 105, -119, -25, -128, 24, 85, -97, 92, 55, 108, -69, -77, -110, 57, -119, -96, 84, -2, -2, 107, 27, -95, 111, 17, -22, -75, -92, 61, -117, 107, -117, 116, 117, -14, 116, 13, -57, -108, -23, 126, -128, 36, -78, -110, -34, -69, -78, -78, 57, 48, -98, -44, 82, -115, 101, -68, -62, -119, 121, -51, 117, -124, -63, 106, -10, -75, -9, 61, -55, 96, 60, -55, 4, 110, -36, 98, -87, 14, -107, 98, -65, -77, -73, -111, -64, -100, -51, 2, -90, -58, 79, -101, -54, -112, -123, 64, -59, -4, -3, 15, -36, -71, 88, 96, -89, -76, 67, -48, 67, 88, -77, -126, -117, -22, -109, -53, 6, -32, 77, 44, 38, 28, 71, 112, 44, 76, 48, 113, -56, -83, 0, 36, -25, -39, 5, 14, 13, -56, 95, -48, -96, -110, -46, -85, -4, -27, -10, -126, 69, -61, 47, -21, 95, -10, -37, 11, -61, -117, -4, 11, -71, 125, -80, 32, -42, 53, -82, 99, 125, -115, -76, -99, -97, 6, -56, 27, 108, 62, 30, 49, -127, -51, -99, 96, 67, -8, -21, -122, 4, 103, 18, 61, 100, 66, -35, -70, -9, 11, -98, -12, 25, -46, 17, 56, 88, 89, -44, 68, 23, 114, -10, 24, -65, 19, -8, -126, -117, 99, -119, 15, 74, 27, -52, 47, -35, 41, 105, 84, -75, -121, -56, 78, -39, 89, 6, -78, 50, 90, 118, -55, 76, -20, 97, -117, 127, -39, -114, -117, -68, -105, 26, -122, 50, 103, 53, -113, 16, 31, 99, 69, 38, -85, 19, -128, -124, -102, -78, 54, 116, -88, 127, 65, 21, 96, 76, 20, -71, 90, 31, -11, 113, -70, -5, 35, -95, -79, 50, 49, 80, 21, -9, -10, 64, -118, -10, 68, -92, 40, -6, -103, 81, -7, 90, -26, -39, 38, 122, 18, 1, 26, -121, -14, 84, 3, -106, 117, 52, 72, 38, 4, -34, -99, 122, -98, -88, -15, 99, -52, -103, -35, -27, 106, 87, -65, -48, -80, 102, -53, 67, -25, 101, 74, 89, 57, -51, 111, 46, -127, 56, -44, 5, -106, -14, 0, -76, 26, 113, -105, 102, -118, -11, -52, 117, -52, 11, -59, -4, -15, 16, -65, 88, -11, -118, 50, -82, -41, 33, 92, -39, -39, -79, 94, -17, 35, -34, 36, -67, -49, 59, -93, -38, -80, -17, -49, -4, 123, 20, 121, -20, -91, -72, -59, 26, -62, 119, 73, 26, 24, 37, 115, 114, 86, 81, -31, -7, -80, -123, 54, -1, 65, 90, 89, 113, -55, -88, -18, -60, 61, -25, 49, 98, 31, 118, -4, 98, 109, -59, -4, 5, 107, -17, -9, 65, -64, 89, -69, -16, 94, 113, 112, 31, 75, 73, 17, -107, 114, 127, -39, 47, -26, -118, 17, -123, -128, -115, 103, 109, -45, -29, -13, -66, 82, 106, 127, -109, 67, -70, 3, 34, -84, -13, -63, 119, -67, 82, -116, -81, 81, -26, 94, -73, -16, -17, -67, -15, -4, -92, -34, 79, 8, 81, -115, -38, 60, -115, -19, -1, -57, 113, -95, -13, -28, -29, -21, 33, -75, -9, 80, -121, 93, 46, -66, -50, -99, -5, 63, 26, 32, -99, -23, -88, 111, -9, 2, 43, 4, 112, -86, 75, 97, -52, -65, -59, 47, 42, 103, 100, -95, 55, 107, 127, -26, -86, -51, 3, 37, -116, -99, -59, -87, 7, -19, -104, 126, 112, 67, 2, 96, 110, -51, 65, -70, 12, -122, 105, -74, 109, 77, -40, 37, 57, -41, -117, 99, 36, 14, 8, 48, 44, 78, 89, -77, -69, 114, -79, -85, 53, 51, -117, 35, -128, 76, 93, 13, 83, 70, 67, 64, 20, -101, -27, -51, -14, -16, -80, -106, 127, 56, 70, 43, 6, 32, 94, 66, 18, -113, 109, -57, 66, 121, 107, 66, 69, 72, -49, 24, 15, -109, -39, -93, -82, 62, -16, 33, -81, 32, 55, -82, -40, -2, 89, 95, -98, 55, 33, 48, 70, 14, 119, 8, 7, 98, -54, -51, 43, 26, 101, -70, 45, -66, -35, 91, 125, 77, -4, -84, -19, -76, -38, 69, 50, -77, 36, 80, 106, -59, 0, 48, 84, -9, -72, -37, -38, 2, 40, -123, -100, 14, -65, 73, 76, 28, 37, 73, -23, -95, 117, 86, -43, -49, 27, -121, 2, -64, 87, -20, 5, -41, -100, -39, 79, -44, 53, -87, 87, -35, -82, 115, 107, -19, 61, 56, -119, -30, 1, -14, 3, -9, -56, 89, 70, 99, 96, -55, -93, 56, 53, 41, -113, 82, -126, 94, -90, 55, -121, 125, -107, -75, 113, -128, 34, 46, 56, 43, -112, -70, -99, 19, 49, -27, -20, -9, -55, -51, 64, -20, -123, -10, -107, -108, -56, -104, 115, -18, 79, 122, -20, 100, -80, -35, 101, 82, -117, 29, -2, -101, 87, 27, 46, 8, -127, -101, -128, -54, -24, 64, 54, -19, -74, 76, 1, -2, 100, -12, 109, 51, -17, -39, 24, 31, 54, -3, -15, 65, -102, 111, 92, 114, 11, 10, -6, 12, 37, -6, 86, -115, -69, 12, -6, -15, -40, 124, 112, -68, -16, 93, 112, 95, -74, 8, -2, 108, -123, 112, 45, -97, 95, 9, -111, -22, -109, 12, 118, 57, -122, 76, 70, -63, -39, -63, 51, 49, -67, 35, 110, 45, 0, 94, 13, 54, -26, -117, 34, -21, 123, -49, 10, 91, 88, 28, -59, 107, -88, -68, 36, -82, -120, -21, -16, -31, 44, -93, -109, 105, 70, -127, 22, -58, 95, -93, 124, -59, -81, 30, 48, -86, 109, -70, -123, 69, 86, -53, 48, 126, 7, -43, -83, 15, 64, 29, 113, -20, 64, -124, -43, 6, -123, 107, 76, 100, -113, 72, -87, -66, -26, 89, -24, -45, -109, -18, -104, 106, 57, 72, 104, -64, -99, -107, 79, 93, 50, 64, -55, -14, 68, 30, 120, 73, 10, 68, 45, 25, 12, 86, 87, 114, 47, -65, -59, 67, 45, -35, 45, -26, -90, 21, 38, -61, 43, -10, -95, -35, -74, -22, 80, 123, -119, 72, 68, 19, 13, -14, -84, -103, -56, -125, -116, 120, -62, -47, 59, 112, 47, -24, -42, 85, 125, 125, -104, 40, -13, -71, -122, 41, 36, 86, 36, 45, 30, -23, -64, -85, 91, -20, -59, -93, -17, -47, -101, 49, 34, 86, 33, -47, -66, 120, -90, -68, 117, -65, 100, -24, -8, 106, -111, -100, 64, 54, 73, -33, -97, -119, 10, 122, -11, 79, -99, 100, -96, -71, 22, 67, -113, -73, -108, -50, -81, -69, 10, -92, -6, -18, 12, 114, -39, 30, -113, -103, -44, 88, -8, -13, 98, -125, -19, -41, 82, 10, -68, 115, 67, 82, 54, 83, -119, 74, -95, -71, -123, 43, -35, -1, -103, 106, -14, -14, 8, 1, 12, 92, -39, -124, -49, -69, -121, 60, 19, 90, -58, 79, 77, -118, 33, 3, 93, 42, -51, 126, 99, -45, 41, -63, 82, 66, -85, -60, -75, 51, 69, 65, 15, -97, 69, 94, -38, 77, 26, 109, 39, 96, 60, -12, 106, -35, 119, 71, -120, -60, 69, 107, 23, -18, -84, -22, -79, -41, 46, -26, -118, -12, -89, 25, 19, 108, -9, 109, 57, -111, 91, -32, 114, 23, 84, 92, 117, 75, 36, 125, -112, -23, 104, 39, 88, -107, -111, -119, -20, 64, -17, -9, -76, 22, -112, 71, 2, 8, 52, -68, 25, 15, 28, 11, -89, -15, -24, -100, -68, -116, -103, -52, -11, -127, 116, -51, -106, -123, -42, 3, 69, 69, 122, 121, -37, -118, 64, 94, 18, -11, -102, -84, -124, 54, 55, -85, -89, -97, -57, -28, -85, -32, 48, 33, -30, 36, 110, -8, 42, -59, 123, -17, -118, 117, -23, -26, -128, -87, -60, 18, 30, -34, 62, 35, -108, -10, 78, -68, 21, -106, 32, 65, -10, -48, -30, 88, 117, -48, -47, 31, 21, -52, -114, 32, -62, -9, -122, -62, 33, -54, 84, -65, 40, 19, 98, 60, -119, 49, 120, 30, 71, 24, -33, -67, 105, 65, -106, 94, -110, -25, -3, 39, 51, 11, -57, 117, -125, -51, -73, 36, 23, -116, 99, -65, 31, 70, 124, 40, -9, 116, -58, -66, 13, 38, -5, -10, -25, 17, -44, -7, 120, 81, -95, 44, -36, -24, 33, -33, 54, 89, -125, -51, 101, 103, 13, 4, 45, 9, -84, -92, -3, -14, -30, -118, -104, 93, 0, 0, -17, 84, 121, -25, 37, -102, -109, -126, 3, 53, -31, -71, 14, -27, 6, -13, -52, -109, 119, 121, 28, -93, -99, -102, 21, -1, -92, 46, -36, 37, -82, 75, -7, -89, -77, -97, -62, -58, -95, 69, 123, 2, 126, 9, 103, 4, 124, -77, 24, 115, -84, -76, -106, -55, -50, 44, 72, -13, -38, -91, -104, 8, 112, 17, 47, -93, 48, 113, -22, 81, 54, -27, -44, 52, 111, -69, -71, 107, -17, 81, 95, 27, -123, 117, 101, -44, 33, 45, 71, 123, 82, 95, 3, 67, -16, -77, 102, -95, -92, -48, 114, 91, 54, -58, 15, 37, 2, 72, 16, 113, 25, -17, 12, 31, -27, -15, 115, -122, -97, 58, -126, 113, 25, 5, 52, -119, 56, 27, -86, 93, 107, -99, 56, 33, -29, -57, -58, 101, -112, 87, 86, 41, -58, -29, -56, 43, 84, -69, 50, 115, 117, 52, 101, 14, -71, 25, 24, 114, -76, 66, 79, -96, 95, 7, 65, -61, 78, -120, -88, 94, 95, 127, 8, -91, -30, 80, 81, -74, -116, 3, -86, -127, -73, -113, 16, -16, 40, -88, -30, 93, 106, -79, 125, 74, 56, 62, -115, 7, 70, -75, -27, 37, -76, 109, 75, 22, 62, 28, 77, 74, -97, 119, 75, -42, -122, -37, 70, 46, 3, -87, 11, -18, -38, 8, -72, -109, -57, -59, 26, -115, -6, 127, 51, 47, 109, -2, -59, 43, -102, -110, -11, -71, -119, -64, 15, -113, 28, -43, 62, -97, -2, -55, 13, 89, 82, 69, 108, -103, -118, 6, -90, 5, 5, 89, -76, -14, -41, -7, -99, -15, 12, 18, 42, 21, 83, -71, 37, -17, 15, -29, 14, -115, 44, -100, 102, -2, 97, 82, 23, 108, -40, 62, -15, 94, 23, 37, -48, 111, -98, -18, -32, 42, -128, -117, -64, 83, -60, 101, -62, 83, -56, 81, 97, 116, 109, 71, -13, 78, 26, -118, 58, 114, 72, -85, 80, -32, 80, -95, -49, 111, 15, 47, 25, 15, 58, 89, -29, 127, 62, 37, 82, -122, -10, 51, 123, -29, -5, -18, -78, -107, -8, 108, -121, -63, -104, 88, 33, 104, 121, 112, 87, 8, 31, -15, -105, -38, -54, -6, -39, -119, -96, -85, -113, 22, 95, -118, 122, -38, -8, -84, -17, 113, -104, -10, -78, -80, -50, 83, -103, -57, 67, 112, 79, -30, -31, 103, 60, 44, -31, -107, 53, 1, -63, 68, -104, -96, 79, -110, -6, -57, -66, 105, -72, -42, -33, -22, 7, 46, -67, 32, 117, -128, 16, 69, -29, 114, 44, -97, 30, -115, -75, -45, 15, -10, -105, 39, 22, 102, 57, -112, -82, 119, 121, -26, -51, -40, 81, 84, -122, -114, -12, 124, -113, -123, 65, -14, 119, -19, 17, 21, -6, 70, 104, -119, -68, 127, 48, 82, 102, -23, 98, -108, -32, 91, -6, 46, -76, -53, 2, -70, -38, 119, -74, -23, 124, 119, 91, 115, -28, -20, 8, 95, -77, -16, 104, -17, -17, 25, -62, -43, -126, -92, -23, -29, -128, 100, -111, -76, -81, 19, -18, 9, 10, 37, 114, 6, 28, 77, -7, -127, -70, -127, 96, -19, -15, 72, 92, 97, -31, -98, -74, -28, -61, 32, 71, -61, 4, 88, -9, 51, -21, 101, -67, 118, 10, -81, -4, -89, 125, 118, -88, -73, 119, -120, 36, -23, 80, 0, -54, -78, 31, 0, 22, 98, -96, -35, -91, 36, -75, 28, -40, 32, 1, 21, 22, -116, 68, -109, -77, 65, -119, -37, 120, -128, -29, 28, -23, -77, -99, 51, -27, 60, -76, 123, 30, -44, -40, 67, 121, 13, -33, -47, -82, 96, 102, 68, 108, 42, 87, -97, -20, 96, -6, -28, 97, 93, -127, -54, -111, -98, 126, -10, 90, -78, -14, -8, 6, 74, -69, -1, -40, 26, 80, 6, -6, 54, -54, -25, -31, -94, 6, 77, -126, -127, -79, 99, 94, -78, -82, 111, -48, -84, -26, -86, -34, 88, 34, 100, 34, 93, -28, 122, -9, -76, 0, 114, 107, 75, -39, -52, 109, 95, -103, 111, 96, -54, 83, 63, -3, -127, 46, 77, -83, -108, 120, 11, 108, 26, -17, 15, -8, 83, 9, 111, -120, -118, 97, 115, 85, -70, -65, 66, -102, -40, 49, 122, 34, 4, 57, -97, 5, -24, 109, 50, -4, 101, -67, -23, -1, 45, 120, 119, 0, 1, 103, 8, 11, 72, -5, -32, -125, 58, -94, -99, -110, 84, -105, 53, -40, 81, 84, 94, -71, 65, 16, 53, 38, 78, -98, -90, -5, -106, -99, 123, 24, -124, 4, -93, 77, 127, 4, 80, 58, 38, 109, 76, -6, -124, 1, 83, 85, -42, 49, -114, -105, -63, 68, 62, -113, 98, 100, 10, 121, -127, 6, 17, -122, -118, 52, 83, -119, -72, 35, 67, 95, 16, 16, -39, 20, -111, -84, -22, -25, 93, -8, -1, -97, -68, -67, -82, -97, -95, 57, -104, -94, -65, 41, -88, -55, -35, 123, -46, 22, 30, -106, -11, -82, 38, 78, 67, 55, 123, -83, -97, 88, 37, 30, 119, 98, 91, -90, -127, 124, 95, -103, -98, -98, 66, -57, -25, -97, -62, 57, 53, 97, 79, -86, -113, -11, 121, 82, -83, 116, 127, -52, 76, 37, 106, 68, 7, 69, 106, 8, 65, 73, 33, 95, 103, -29, -90, -50, 2, -23, -121, -72, -54, 87, -30, -39, -52, -37, -84, -7, -49, -85, 69, -100, 80, 47, 96, -41, -12, 74, 95, -75, 19, 0, -107, -6, 99, -69, 72, -26, 36, 79, 30, 110, 38, -128, -56, 115, -36, -12, -20, 43, 31, -78, 71, -16, 97, 39, 71, -42, -15, 39, 11, -124, -89, 32, -2, -117, 92, -58, -15, 0, -106, -113, -17, 60, -113, 55, 47, -21, -85, -100, -105, 74, -50, 94, -70, -81, 6, -126, 5, 119, 41, -111, 124, 80, 49, -6, 91, 13, 65, -52, -114, 87, -37, -3, 19, -21, -76, -61, 86, -33, -33, 109, -87, 45, 76, -28, 92, -46, -26, -30, -55, -113, -13, -59, 95, -92, 64, 59, 50, 1, -121, 64, -40, -29, -67, 107, 78, -15, -82, 36, 80, 13, 18, 121, -70, -34, -35, -105, 48, 67, -7, 121, 82, 108, -65, 50, -112, 127, -19, 66, 0, -12, 2, 88, 87, 63, 67, 37, -80, 114, -54, -128, -1, 92, 122, 58, -70, -41, 81, 106, -101, -54, 99, 109, -74, -94, 31, -58, -95, -116, -119, 33, 1, 11, -7, -40, -53, -67, 126, -5, -81, -56, -4, 46, -92, -10, -24, -34, 77, -71, -56, 104, 3, -85, 86, 57, -50, -11, -128, -17, 2, -119, -111, -125, 20, 10, -37, 95, 71, -39, -37, 118, 33, 87, 37, 69, -51, -115, -93, -102, -57, -21, -125, 74, 23, 89, 4, 101, -50, 4, -44, 80, 13, -27, 83, -95, 112, -81, -127, 55, 8, -36, 46, -86, -77, -45, 111, 0, -32, -109, 26, 39, -2, 29, -14, -107, -10, 118, 122, 69, -6, -49, 21, -121, 52, -23, -88, 36, 24, -87, -36, -96, 5, -118, -54, 56, -35, -70, -72, 61, -51, 83, -27, 75, -16, 87, 97, 103, 77, 91, 44, -57, -86, -63, -50, 95, 42, -10, 3, -62, 32, 95, -29, -91, 105, 45, 94, -58, 103, -106, -124, -76, 105, -23, -128, -38, -64, 97, -63, -115, 60, 109, -44, 103, -82, 34, 70, 89, -104, -55, -101, 56, -87, -2, 94, -110, -84, 60, -39, -109, 82, -35, -56, 60, 70, -56, -106, -122, -87, -41, -109, 101, -60, -25, 76, -14, -119, 18, -53, -95, 92, -25, 90, -123, 101, 56, -105, -111, -12, -16, -91, -58, 77, -19, -126, 19, 53, -104, 25, 94, -17, 44, 67, 51, -109, 16, -90, -100, -94, -15, -66, 126, 88, -104, -125, 62, 80, -101, 79, -60, 11, 116, 10, -39, -31, 13, 108, -106, 37, 6, 116, -107, -78, 56, 72, -58, -56, 110, -30, -22, -32, 32, -23, -72, 56, -20, 118, 8, 7, 70, 76, -109, 58, -41, -20, -100, 100, -40, -78, 9, 94, -89, 30, -111, 95, -25, -41, -89, -43, 57, 17, 53, -38, 122, 110, -110, -25, 100, 27, 110, 42, -25, -127, -27, 62, -19, 1, 34, 70, 51, -84, 36, 90, 74, 53, 57, -79, -116, 96, 7, 70, -14, -68, -96, -20, -86, -78, 83, -113, 77, 66, 57, -75, 67, -98, 115, -79, 31, 22, 119, -45, 66, 27, -83, 12, -47, 103, 62, -35, 71, -59, -93, -71, 1, -61, 38, 44, -10, -7, 59, -61, -69, -12, -8, 127, 19, -20, -80, -78, -126, -89, 5, 68, 66, 51, -48, -109, 26, -114, -15, -31, -45, 20, 27, 85, 88, -63, 1, -50, 58, -68, 17, 118, 48, -118, 117, -61, -10, -91, -10, -8, -52, 123, -68, -114, 46, 12, -94, -56, 27, 19, 42, 110, -89, -59, 67, 127, 6, -60, -51, -64, 0, 95, -74, -79, 105, -85, -12, -33, -48, 106, 87, 28, 102, -109, 43, 20, 31, 77, 93, -70, -32, 7, -87, 7, 76, 108, 7, -46, -79, 84, 18, 49, 51, 73, 98, 28, 116, -41, 123, -59, -63, 82, 97, -89, 101, 12, 60, 5, -39, 25, 63, 57, -96, 104, -63, 108, 85, 72, -66, -122, 28, 80, 55, -48, 25, 26, 108, 14, 113, 104, 83, -78, 58, 52, -38, 32, -63, -106, -91, 26, 47, 100, -44, 79, 77, 21, 59, 34, -35, 121, 40, 121, 73, -33, -55, -29, 121, -74, 113, 106, -98, 68, -99, 88, -8, -9, -8, 57, 13, 29, -44, -68, 2, 40, -117, -49, -67, 70, 113, 26, 63, 25, 19, 8, 120, 93, 107, 114, -109, 92, 92, -79, 32, 121, -119, -103, -16, 2, 82, 125, -97, -90, -71, 33, 78, -60, 112, -117, -118, 97, 37, 73, -6, -71, -46, -13, -106, -67, -27, -87, -102, -63, -38, 58, -69, -29, 83, 43, 101, 38, 41, -123, 76, 98, 38, 27, -89, 23, 38, -79, -8, -52, 123, 115, 5, -51, -26, 27, 10, 75, 68, 36, -116, -98, -33, -57, 1, -78, 115, -25, 88, 28, -20, 37, -2, -110, -64, 37, 41, 102, 87, -94, -78, 82, -107, 55, -97, -5, -46, 41, -58, -106, -50, -46, -76, 45, 26, 54, 95, 13, -99, 56, -87, 9, -35, 39, 27, 29, -51, -59, 3, -92, -25, 54, 118, -4, -19, -107, 119, 64, 62, -67, 86, -116, 15, -117, 57, -87, 65, 25, 54, 94, -47, 95, -25, 46, 7, -126, -53, 84, -57, 78, 120, 46, 4, 110, -86, 114, -125, -95, 50, 65, -34, 8, 78, 110, 19, 7, -105, -44, -96, 78, -78, -15, 45, 25, -97, -76, 28, -22, -120, 99, -71, -128, 18, 61, 110, 60, 47, 113, 94, -31, 51, -68, 106, 1, -86, -3, -120, -62, 82, -87, -112, -124, 26, 61, 30, 58, 114, -70, -92, 122, -99, -35, 123, 47, -101, 105, -20, 74, 91, -54, -84, 14, 6, -106, -113, 49, 19, -105, 115, -27, -64, -125, -22, 91, 64, -120, 21, 50, -62, 57, 45, -33, -105, 40, -113, -78, 17, -5, 124, -20, 69, -88, 122, -53, -66, -119, 124, 82, -95, 111, -73, -31, 114, 33, -68, 51, 41, 81, -27, 107, 11, -110, -53, 34, 58, -38, 84, -52, 85, 80, 56, 26, 121, 51, 101, -73, 60, 98, -119, 93, 81, -63, -65, 68, 98, -5, -9, 12, -51, 92, -9, 88, 111, 66, -6, 41, -100, -50, 117, 113, -98, 46, 11, -105, -31, -15, -49, -99, -45, -40, 123, -92, 25, -70, 104, -4, 53, -33, -120, -126, -68, -1, 90, -85, -62, -44, 84, -34, 34, 74, -48, 65, -8, 91, 88, 89, -52, -89, 118, 31, 0, 113, 68, -103, -85, 44, 21, 97, -116, 29, 99, -56, -99, 62, -13, -33, -110, -57, 61, 53, -111, -115, -10, 9, 105, -50, -30, -75, -10, -39, 85, 118, -54, 25, -113, -10, -59, 37, -41, -47, -62, -70, 25, -33, 120, -116, 62, -117, -44, -4, 64, -27, 9, -74, 111, -14, 4, -47, 40, 122, 42, -3, 112, 117, -106, -128, -21, -37, 37, 66, 45, 103, 124, -58, -57, 117, -45, -123, -128, 39, 1, 64, -116, -117, 118, 123, -3, -6, -51, -91, -11, 119, 34, -27, 108, 56, -27, -41, -108, -118, -103, 65, 114, -106, -121, -71, -117, -38, -66, -117, -127, 64, 75, -114, 75, 65, -119, -56, -69, -42, -18, 48, -50, -112, -106, -70, 73, -5, 18, 93, 6, 43, 30, -8, 65, 37, 49, 76, -128, 111, 87, -127, 47, 34, -113, -6, -29, -103, 67, 31, -17, -79, -49, 61, -63, -27, 120, -118, 97, 10, 103, -25, -75, 5, 95, 119, -85, 16, 67, -85, -1, 27, -84, -81, -67, -68, 41, 33, -43, -20, -64, 68, 29, 15, 2, 95, 117, -6, 105, 86, -124, 81, -67, -71, -42, -100, -80, 1, 44, 116, 44, -85, 15, 89, -38, 76, -107, -124, -19, -22, -16, 45, -82, -114, -67, 48, 109, -78, -86, 86, -120, -82, 39, -59, -24, 126, -31, 24, -1, -115, 12, -84, -72, -101, -123, 19, 104, -102, 23, -43, 4, -121, -125, 50, -107, -64, -29, -126, -14, 13, 89, -6, 60, 0, 63, -92, -2, -96, 60, 126, -83, -55, -86, -27, -28, -81, 120, -52, -55, 15, 34, 77, 23, 37, -1, 44, 101, 98, 47, -41, -16, 8, 81, -84, -120, 16, -48, 7, 48, -116, 5, 93, -43, 47, -62, 58, 94, -69, -122, -89, 74, 40, 116, -31, -51, -13, -114, -78, -42, 61, 9, 70, -59, -38, 114, -51, 106, -62, 84, 26, -50, -39, -9, 36, -120, 58, -34, 102, 117, -28, -115, 63, -115, -127, -95, -38, -11, -81, 13, 75, 108, -106, 17, -79, -15, 3, -2, -37, 69, -45, 118, -109, 44, -19, 55, 53, -89, -107, 27, -100, -6, 41, 92, 7, 42, 125, 97, -97, -84, -18, 106, -104, 5, -5, -55, 118, 126, 71, -47, 67, -102, -57, 87, 71, 53, 14, -4, 92, 36, -105, 121, -98, 64, 85, 37, -21, 82, 6, 10, 126, 117, -11, -106, -6, 112, -33, -16, 111, -90, 65, 50, -63, -119, 9, -120, 62, -104, 4, 26, 60, 27, 19, 90, -36, -24, -1, 71, -70, -123, -47, -72, 122, 70, -50, -12, 55, 45, 100, 38, 84, 38, -40, -107, 47, 98, -99, -19, 122, 33, -121, 54, -68, 27, 16, 24, -125, -113, -33, -66, -108, 49, -10, -113, -9, 69, 3, -82, -14, -24, 84, -58, -114, -83, -37, 61, -113, -8, -86, -119, -103, -79, 63, -42, 76, -49, 110, 80, -34, -50, -114, -14, 127, 4, 1, -10, -55, -123, 37, 60, -19, -7, -126, -5, 38, -34, -72, 53, 86, -30, 62, 112, 19, -3, -58, -32, 76, -76, -80, -86, 2, -66, 29, 1, 66, -98, 120, -116, -93, 29, 72, 16, -106, 74, -117, 61, -88, -61, -14, 127, 37, -79, 111, -71, 46, -75, 25, -5, -23, 73, 37, 108, -121, -62, -19, 73, -31, -27, 85, 4, -126, 29, -107, -103, -24, -96, 86, 16, -28, -56, 15, -119, -7, -2, -62, -88, 51, 91, 35, -99, 36, -56, -119, 43, 11, -10, -11, 108, 92, -54, -16, 94, 104, 5, 119, -48, 38, 77, 96, -118, -106, -16, -109, 15, 110, -42, 55, 34, -79, -38, 63, 86, 35, 72, 1, -82, -66, 118, -102, -102, -63, 10, 121, -87, -112, 112, -7, 54, 62, -39, 64, 84, 73, 83, -29, 56, -87, -101, -38, -37, -11, -103, -79, -104, 97, 50, -58, -97, 41, -32, -70, 106, 107, -77, -109, 123, -93, 12, 49, 97, 101, -15, 53, 47, -60, -103, -25, -18, -76, 65, 73, 41, 90, 122, 66, 59, 44, -120, 90, -43, -23, -108, -65, -44, -57, -46, -49, -21, 94, -128, -52, 68, -15, -126, -13, 53, -101, 90, -93, -49, 27, 108, 120, -11, 102, 58, -80, 19, 67, -118, 104, -84, -97, -88, 0, -26, -6, 79, 81, -39, 79, -98, -99, -64, -96, 16, 117, -69, -22, -103, 10, -123, -123, 2, -6, 108, -67, 42, -1, -128, 52, -25, -84, 83, 15, 44, -70, -118, -5, -117, -29, -54, -87, 0, 10, -55, -112, -1, 4, -6, 24, -114, -1, 30, 17, 121, 10, 78, 35, -119, 78, -41, -16, 122, -85, -128, 38, -27, -118, -95, -16, -19, -21, 26, 109, 117, 99, 125, -12, -24, -9, -115, -10, 118, 43, -121, 111, -75, 85, 18, -66, 35, 105, 46, 29, -108, 46, -61, -7, 56, -28, 106, -91, 79, 4, -110, 68, -25, -113, -71, 79, 6, -58, -58, -4, 113, -51, -21, -90, -93, 125, -28, 70, 103, -110, -28, 123, 65, 39, -11, -7, -116, -33, 31, 91, 99, 49, 32, -54, 65, 89, -102, -57, -97, -32, 68, -112, 45, -81, -74, 80, -83, 26, 23, -108, 44, 123, -113, -19, 34, 4, 103, 46, 99, 6, 10, 70, -73, -86, -111, 120, -125, -85, -64, -94, 11, -124, -78, -72, -77, -24, -119, -32, -126, 32, -12, 46, 27, 4, -100, -67, -120, -125, 108, 108, 9, -10, 50, 64, 32, 67, 57, 35, 110, 121, 69, -7, 125, 119, 50, -80, -33, 59, 17, -31, -37, -123, -113, 118, 9, -85, -77, 18, -82, -97, -2, 55, 21, -80, -8, -75, 116, -79, 88, 98, -86, 29, -36, -89, 20, -114, -41, 115, 73, 104, -44, -92, 110, -28, -102, -9, 15, -51, -119, 62, -19, 7, -11, -126, 56, 109, -72, 44, -98, -112, 14, -56, 46, 106, -17, -62, 120, 71, -74, 65, 47, 10, 101, 29, 110, 127, -107, -2, -51, -98, -68, 58, 38, 49, 60, -34, 31, 116, -118, 61, -123, 24, -122, 51, 3, -11, 117, -5, -68, -85, -67, 108, 54, -94, 9, 36, -94, 30, -94, -17, 61, -34, -87, -29, -112, 101, 65, 47, 90, 75, -20, 95, -29, -14, 18, 102, 104, 7, -30, -92, 51, 31, -112, -23, 65, 26, -115, 99, -72, -80, -46, 117, 14, -5, -40, 30, -31, -103, -51, -69, 100, 58, -102, -56, -84, 44, -82, -108, -77, 16, -71, 102, -81, -55, -49, 113, 99, -35, 84, -100, 13, -89, -111, -101, 34, -22, 58, -125, 3, -121, -66, -24, 65, -40, 48, 110, -124, 94, -126, -72, -17, -69, -98, 30, 5, -18, 15, -24, 75, -28, 4, -40, 11, 22, -13, -83, -128, -83, -79, 3, -75, -17, 107, 118, 72, 27, 100, 76, -6, 103, -124, 105, -94, -93, 7, 39, 17, -105, -112, -36, -5, 20, 52, -122, -86, -89, -77, -86, -43, -28, 46, 10, 84, 25, 0, 28, -75, -27, -24, 47, -52, -19, 24, -18, 16, -97, -106, -95, -74, -90, -3, 49, 58, -79, 55, 101, -40, 107, -113, 45, -49, 61, -73, -93, -41, 56, 63, 12, -99, -88, -69, -23, 21, 83, 87, -91, 114, 109, -58, -87, -109, 67, 90, 78, 116, 18, 51, -52, -3, 66, 122, 76, 0, -79, 112, 87, 105, 47, -29, -122, 87, 30, -17, -20, -15, -57, 17, -29, -76, 87, 12, -56, 26, -25, -106, 14, 121, 73, 91, -10, 11, 85, -62, -117, -122, -78, 98, 112, 98, -59, 118, 57, 99, -26, -90, -44, 45, 55, 56, 97, 15, -60, -87, -87, 43, -65, 56, 36, -120, 19, -102, 20, -24, -35, 31, -18, 15, 2, -34, -15, 71, -43, -85, 43, 59, -47, 127, -24, -120, 55, -55, 23, 124, -13, 65, 39, 50, -7, -52, 59, -116, -26, -49, -12, 67, 110, 98, -45, -16, -63, 68, -72, 22, 111, 99, -47, -64, 98, 57, -55, 26, -126, 96, 22, -11, 33, -67, -88, -102, 9, 99, -90, 112, -78, 26, 51, -96, -3, -122, 17, 62, 75, 73, -44, 58, 44, 37, 123, 14, -34, -60, -88, -32, -92, 62, 86, 70, 124, 126, 96, 5, 97, -121, -11, -109, 33, -87, -77, -98, -81, 68, 92, 122, 13, -80, 53, -71, 85, 48, 72, -77, 116, 112, 20, -104, 47, -22, 94, 43, -24, 63, -80, -55, 70, 38, -36, -25, 79, 15, 6, 126, -44, -30, 121, 97, 19, 46, -101, -24, -34, 99, 28, -46, 83, -80, -22, 2, 26, -55, -83, -126, -120, -34, -53, 78, -124, 39, -75, 83, -74, 59, 81, 10, -98, 74, -20, 49, -8, 7, -103, 86, -22, 53, -88, -67, 101, 19, 64, -1, 92, 109, 1, 100, -53, 76, 50, -49, -13, 103, -94, 42, 35, 116, -76, 65, 62, 32, -14, -73, -89, 11, -115, 17, -63, -74, 79, -90, 73, 15, 38, 37, -4, -89, 9, 72, 116, -69, -105, -25, -94, -70, -111, 69, -82, -58, 6, 108, 102, 120, -93, -114, 4, -79, 31, 69, -25, -18, 107, -80, 125, 17, 85, -6, 57, -34, -62, 45, 25, -39, -108, 59, 19, -90, 1, 65, -20, -121, 46, -46, -128, 81, -32, 4, -126, -128, -55, -23, -18, -76, 25, -20, 70, -18, 102, -1, 76, -88, -84, -27, 1, -64, -95, -107, -26, 34, 86, 82, 41, 4, -91, 41, -42, 5, -83, -40, 5, -10, 66, 116, 43, -37, -32, -15, 74, -58, 112, 22, -18, -100, 124, 111, -36, -99, -124, 67, 63, 91, 21, -24, -33, 58, -110, 53, -64, -65, -114, 69, 54, 80, 57, -31, -85, -103, 82, 117, -33, 66, 12, 77, 94, 8, 61, -70, 37, 65, 125, -28, 28, 19, 76, 124, -51, 94, 49, 13, -98, 63, -45, 84, 15, -116, -75, 59, -90, -121, 48, 5, 73, -68, -45, 39, 68, -112, 97, -23, 81, 95, 77, -18, -14, 26, -22, 63, -8, -101, -51, 22, 91, 32, -22, -22, 44, 31, -91, 82, 38, 86, -40, -17, -110, 43, -106, 87, 59, 120, -64, 12, 87, -114, 122, -55, 40, -28, -120, -96, 0, -43, 55, -37, 117, -95, 69, 34, 65, 107, -12, -25, 65, 76, 87, 83, -9, 109, 42, -78, 101, 107, 63, 60, 121, 57, -123, 33, -98, -114, 65, 30, -29, -8, 121, -39, 26, 62, 123, -37, 41, -17, 66, -22, -68, 25, -66, 51, 7, 104, 102, -20, 83, 37, -87, 76, -34, -82, -19, -4, -68, -81, -102, 32, 39, -109, 121, -63, 82, 116, 28, -5, -29, -33, 102, 31, 120, -92, -45, -1, -116, -71, 108, 96, 94, -107, 44, -68, -61, -102, 57, 0, -55, 83, -96, 112, 103, -103, -78, 57, -115, 78, -76, -16, -83, -102, -112, -90, -66, -29, 37, -53, 28, 17, -85, -6, 38, 87, 54, 106, 113, -17, -22, -70, -61, 10, -85, -86, 35, -35, 99, 48, -85, -105, -96, -39, -78, -80, -1, -16, 19, -92, 59, -81, 54, 102, 41, -36, 62, -32, -58, 47, 79, 48, 106, -110, -70, -107, -68, 93, -14, -97, 13, 29, -73, 46, 118, -23, 94, -11, 89, -14, 26, 21, 33, -48, -5, -53, 44, -71, 43, 115, 105, -6, 35, 83, 13, 94, 104, 73, 59, -38, 105, -55, 119, -96, 119, 110, 9, 85, -29, -30, -57, 125, 119, 105, -51, -13, -76, 122, 44, 95, 109, 21, -39, 16, -24, 102, -18, -48, 48, -86, 42, 25, -13, 34, 57, -22, 16, -62, -65, 115, 36, 7, 113, 28, -16, -66, -113, 36, -72, 59, 3, -91, -47, 92, 54, 57, 67, -92, -118, -13, -50, 52, -116, 65, -42, 69, -85, 102, -121, -21, 90, 43, 114, 75, -57, -30, -119, -42, -122, -62, -110, 9, -25, -29, -27, -99, -100, -88, -62, -90, 27, 16, 91, 39, -46, -79, -20, -3, -104, -13, 104, 114, -97, 90, 61, -26, -68, 70, 61, -62, -120, 79, 75, -16, -78, -79, 13, -50, -39, 79, -11, 117, -32, -48, 28, 50, 1, -119, -81, 25, -4, -104, 11, 27, 114, -56, -126, -81, -113, 63, -15, -105, 14, -67, 7, 64, -18, -107, -114, 71, 100, 3, 60, -60, 83, -39, 118, -43, -30, -90, 110, 94, -66, -6, -6, -80, 66, -4, -33, 81, -69, 81, 105, 73, -114, -16, 9, -4, 5, 23, -61, -22, -101, -128, 46, 110, -39, 37, -61, 59, 75, -78, 25, -119, 44, -109, -71, -18, 15, 25, -64, 74, -22, -87, 19, -8, 25, -100, 116, -97, 52, -73, 9, 79, -73, -73, 61, 16, 92, -127, -53, 39, -77, 101, 48, 95, 120, 106, -51, 8, 3, 13, -46, 109, 54, 102, -27, -48, -126, -39, -17, 54, 16, 120, 5, 72, -81, -61, -40, -116, -60, 36, 51, -9, 9, -28, -42, 1, -50, 35, -119, 81, -79, -36, 62, 103, -62, -93, -73, -60, -4, 38, 123, -116, 30, 0, 84, 78, 67, -83, 90, -121, 81, 13, -2, -38, 113, 84, 91, -65, -8, 101, -112, 41, -63, 78, 16, 3, 113, 72, 71, -19, -18, 66, -6, -115, -61, -50, 91, -122, -5, 53, -114, -52, -62, 12, 38, -76, -31, 2, -13, 89, -25, 4, 2, 40, -46, -110, -85, -60, 90, 114, 49, -55, 53, -85, -42, 120, -6, -79, 126, 117, 102, -116, -62, -88, 25, 104, -36, 122, -22, 80, 83, 81, -44, -43, -7, 38, -25, 36, 106, -62, 23, 28, 11, -52, 71, 97, -60, -63, -110, -62, -73, 120, -49, -7, -96, 104, -31, -3, 98, 76, -51, 53, 29, 33, -118, -105, -57, -15, 59, -78, 51, -46, 78, -66, 30, 21, -97, 98, 87, -79, -91, -114, -87, -12, 7, -54, -36, 104, 71, -66, 52, -108, 115, -46, 53, 125, -23, 124, -18, -92, -82, -94, -9, 124, -32, -107, 18, 0, 120, -23, 49, -99, -9, 91, 17, 126, -91, 109, 102, 108, -85, 27, -128, -98, 109, 53, -101, -42, 49, 9, -6, 96, 43, 113, 92, -116, -121, -18, 12, 127, 87, -67, -100, -50, -104, 45, -52, -67, 26, -77, -87, 69, 78, -87, 99, 59, 94, 126, -111, 16, 7, 11, -16, -77, -3, -52, -65, 4, 59, 75, 3, 18, -120, 31, 97, -95, -52, -83, -34, 102, -32, 8, 43, -82, 49, 14, 105, 16, 12, 122, -96, -109, 6, 16, -58, -125, 92, 5, 7, 23, -48, -118, -86, -39, 41, -117, -6, 117, -72, 88, 91, 25, -32, 6, 71, -110, -108, 49, 34, 32, 43, 66, 51, -79, -46, 122, -76, -82, -1, 59, 70, 80, 69, 112, -87, -18, 123, 35, -29, -77, -5, -66, 76, 92, 68, 20, 110, 88, -59, 16, -8, 112, -46, -84, -94, 36, -90, -42, 82, 37, -110, 24, -11, 87, 8, 30, -58, 3, -63, 41, 55, 61, 104, 3, 25, 44, -105, 7, 5, -36, -105, 125, -51, -23, -87, -17, -115, -49, 69, 95, 117, 87, -8, -22, 47, -128, -119, 117, 4, -54, 30, -69, -121, 6, 62, 32, -77, 86, -89, 56, -78, -66, 53, -1, 39, 95, 110, 52, -82, 52, 20, -93, 11, -116, 14, -70, -116, 23, -81, 16, 97, 78, 75, 105, -44, 10, 9, 7, -32, 49, -65, 18, 111, 117, -110, 23, 84, -128, -53, -126, 52, 95, -90, -64, 107, 52, -6, 120, -53, 42, 8, -84, -8, -44, -107, 76, 94, 31, -44, -66, -48, 19, 80, -65, 8, 98, 86, -36, 99, -94, -33, 23, -127, 5, 87, 109, -71, -46, 101, 4, 124, -19, 48, -12, 65, 70, -64, 31, -27, 20, 93, 53, -88, 46, 116, 48, 16, 75, -115, -13, 109, -20, -117, 110, 113, 98, 91, -86, -76, 64, 46, -80, -82, -34, 36, 111, -92, 101, 15, 9, -7, -20, -66, 33, -102, -77, -46, 43, 126, -33, -98, 107, 75, -87, 89, 60, -116, 53, 102, -64, -11, 20, -15, 35, 114, -107, 19, -105, 122, -94, 32, -12, 14, 95, -107, 41, -110, -25, -44, -112, 70, -14, 123, 17, 28, 84, -51, 40, 9, -77, 104, 127, 71, -39, 34, 58, -17, -75, 81, -23, -41, -15, 93, 102, -48, 115, 15, -30, -38, 99, -14, -95, -43, -19, 50, 113, -62, -128, 25, 75, -77, 2, 74, 123, 91, -19, 53, -54, 34, 6, 52, 122, 119, 17, 96, -56, 4, -17, 42, 95, -46, -99, -128, 39, 10, 50, 25, 76, 50, -78, 24, 102, 52, -30, 97, 16, 79, 22, 90, -14, -100, 14, -20, -109, -96, -52, -37, 36, 59, -122, 3, -115, -93, 3, 52, 45, -74, -51, -6, 104, 0, -110, 78, -76, -12, 47, 68, -60, -59, 31, 54, -31, -83, -94, -11, -51, -18, 80, 114, -87, 86, -11, -74, 121, 121, 106, 39, -81, -72, -95, -105, 56, -77, 102, 108, 39, 21, 49, 107, 91, -48, 33, -68, -3, 67, 49, 75, -79, 2, 61, -38, -40, -78, 16, -46, -85, -5, 121, -38, 51, -102, -14, -21, -51, -40, -41, 116, 109, -120, 96, 72, -40, 1, -123, 86, -59, 54, 33, -10, -72, -34, 81, 17, 16, -31, 99, 60, 92, 92, -106, 15, 118, 8, 122, -61, 96, -46, -73, 78, -38, -105, 22, 51, 25, 27, 9, 94, -46, -86, -44, 10, 8, -91, -101, -104, 7, 126, 84, -29, 90, 107, 115, 80, -13, 109, -109, -44, -65, -53, -94, 26, -30, 56, -51, 123, -44, 86, 89, 38, -128, -82, -80, 8, -45, -52, 32, 90, -54, -11, -66, -91, -32, -79, 117, 83, -98, -119, -89, -34, -44, -55, 120, 54, -126, -59, 50, -42, -101, 11, 124, -101, 57, -84, 35, -115, -8, -61, 103, 67, 56, -91, 104, -104, -42, 93, 108, -11, 102, -109, 83, -70, -35, 75, 113, -33, -112, 35, 53, -85, -82, 49, -58, 104, 93, 105, 117, -42, -84, 92, -103, 101, -126, -127, 125, -40, 94, 105, 77, 69, 125, 32, 127, -38, -21, 112, 57, -5, 19, -18, 38, 66, -97, 108, 42, 124, 85, 31, -46, -126, -5, -21, 103, -3, -20, 100, 86, -53, 78, 35, -112, 75, -60, -113, -91, 47, -128, 94, -85, 19, -52, 81, -43, -21, 62, 127, -25, 19, 30, 58, 21, -102, -91, -4, 23, 18, -31, -19, 93, -81, -111, 109, 122, -43, 124, -97, -124, 124, 125, -81, 16, -55, -127, 101, 52, 63, 101, -101, -46, 3, 85, 104, 29, 123, -28, -75, 13, 69, 34, -22, 116, 51, -41, 110, -120, -45, -115, -115, -48, -118, -68, 96, -45, -67, 69, -121, 124, 42, -93, -49, -82, 120, -73, 75, 115, 27, -128, 0, -31, 35, 106, -43, -42, -63, -60, -33, 21, -47, -20, 101, -36, 40, 69, 47, 102, 10, 55, 98, -75, 90, -79, -29, 82, -24, -82, 70, -124, -81, -58, -27, 82, -79, 58, -88, -14, 126, 7, -121, -48, 115, 108, 44, 28, 49, -37, 2, -68, -110, -28, -15, 108, 22, 84, 63, 126, -126, 5, -126, -79, 75, -25, -125, 124, -94, -84, -17, -96, 51, -10, -16, 39, -29, -100, -61, -108, -8, 69, -48, 10, -87, 65, -9, 63, 21, -74, 62, 24, 59, 64, 73, 6, -88, 77, 3, -54, 121, 114, -22, 44, -24, 91, -45, 75, 119, 22, 96, -17, -37, -80, 122, 5, 114, -15, -60, 7, 39, -126, -97, -30, 67, 105, 104, 107, 54, -21, -75, 47, -35, 31, -37, 70, -6, 47, 17, -14, -59, -15, 97, 33, 34, 91, -90, 20, -52, -22, -101, 115, -19, -69, -43, -80, -92, -66, -101, 90, 41, -48, 9, -121, 111, 100, 77, -22, 19, -34, 92, 89, 80, 61, -6, -14, 25, 32, -122, 101, -118, -95, 89, -9, -36, -82, 39, 0, -20, 66, -38, -106, -110, 99, -99, -126, 72, 106, -20, -37, -56, -56, -76, -104, -123, 46, 10, 30, -50, 16, 4, -39, 50, -35, 80, -114, 11, -8, 15, 120, -70, 105, -114, -51, 77, -85, -49, 21, -107, 59, 112, -35, -125, -91, -10, -120, 83, -128, 39, -94, 17, -85, -5, -61, 8, -53, -47, -109, 67, 96, -117, 126, 74, -103, -53, 23, -60, 26, -84, -39, -43, -100, 55, -40, -63, -83, -32, -107, -83, -121, -73, 62, -78, 50, -127, 58, 125, -45, 78, 65, -77, 89, 63, 125, 115, -118, 20, -73, 36, 64, 17, 121, 93, -56, -47, -98, -11, 49, -77, 34, 57, -22, -31, 107, -100, -30, 38, -102, 53, -12, 91, 105, -51, 26, 102, -64, 36, -5, -8, -56, -69, -119, -63, -104, -47, 18, -73, 70, -61, -22, -24, 124, 85, 73, 104, 113, -84, 14, -117, 97, -126, 102, 74, -49, 0, 49, 16, -92, -84, -120, -20, -25, -111, 45, 0, -30, -65, 55, -88, 3, -95, 16, -1, 118, -38, -25, 104, 6, 117, 115, -25, 119, 90, -78, -57, -38, 99, 87, -1, -113, 95, 107, -10, 112, 25, 118, -46, 88, 45, -6, -37, 79, -118, 91, 69, -28, -62, 45, 106, -72, 33, -46, -81, -5, 4, -10, 85, -25, -51, -44, -10, -84, -64, 108, -100, 89, 99, -18, 49, 16, 104, -115, -33, 115, 104, -91, -41, -86, 82, -62, -30, -13, 20, 18, 110, -104, -120, 68, -1, -42, -104, 117, 2, -40, 97, 31, -79, 68, -115, 99, -43, 118, 112, 52, 105, 88, 89, -64, -126, 44, 2, -27, -97, -106, 119, -114, -82, 127, 82, 45, -43, 106, 34, 88, -61, 4, -9, -12, -56, 4, -41, 29, -6, -57, -46, -29, -97, -85, 36, -94, 87, -90, 7, 119, -67, -2, -123, -21, -3, 87, -103, 83, 65, 59, 43, -124, -65, -94, -7, 8, 38, 80, -91, -95, -104, -9, 4, -73, 35, -88, -39, -6, -49, 96, -15, 12, -34, -10, 119, 92, -51, -112, 47, -113, 76, -38, -109, -117, -4, 12, 19, -94, -35, 57, -61, -11, -80, 72, 44, 83, 112, -122, -50, -65, 102, 63, 75, -59, -74, 67, -95, 3, 83, 80, 18, 31, -86, 38, 43, 38, -78, -66, 72, 15, 119, -116, -124, -88, 84, 49, 123, 68, 55, -55, -124, 29, -119, 79, 98, -65, 18, -125, 66, -26, 83, -43, -123, 125, 123, 48, 35, -83, 111, -20, 61, 102, -8, 65, -114, -52, -14, -118, -112, -87, -45, -108, 71, -36, 100, 41, 27, -10, 45, -34, 92, 0, 51, 98, -2, 46, 18, -95, 91, 1, 13, 24, -24, -123, -38, -10, -47, 76, 0, -30, 118, 84, -10, 61, -80, -38, -26, 76, 81, -109, -86, 45, 20, 93, 15, -110, 11, -94, -77, -26, 35, 65, 127, -117, 70, -39, 2, -104, -91, -126, -6, -101, 86, 112, 88, -121, -53, -65, 83, -100, -46, 125, 73, 102, 90, -39, 120, -27, -5, -84, 75, -98, 109, 74, -86, 51, -93, 44, 75, -55, 46, -59, -28, 5, -74, -67, 12, 1, -4, -33, 29, 78, -36, -26, 53, -74, 63, 45, 27, -70, 89, -26, -39, 70, -79, 3, -6, -44, -81, -59, 29, 93, 11, -126, -30, 65, -65, 110, -62, 59, -51, 95, 9, 41, -59, -66, 95, -123, 108, -6, -65, 69, 97, 24, 12, -110, -101, -122, -26, -54, -53, -124, -88, 86, -122, 10, 23, -59, -7, 89, -128, 70, 56, 9, -16, 126, 72, -49, -125, 52, 74, -62, -7, 43, 91, -123, 61, 118, -117, -93, -63, -41, -89, -23, -83, -83, 115, 69, -14, -20, 30, -14, -77, -41, 124, 35, -43, 68, 114, -40, -8, 60, 26, 113, -25, -11, 119, -92, -20, -126, -56, 45, -39, -17, -106, 7, 29, -119, -52, -113, -10, 106, 2, 41, -63, -2, -52, 22, -62, -66, 110, 58, 123, 9, 43, -30, 126, 34, 7, -22, 37, 79, -105, 126, -66, -83, 5, 91, -73, 81, 107, 45, 60, -19, -42, 125, 107, 34, 20, -83, 96, 2, 103, 91, -117, 18, -66, -118, -75, 69, -12, 90, 20, 12, 88, 82, 57, -34, 46, 112, -81, 25, 29, 107, -122, 115, 105, 113, 21, -3, -98, -10, 127, -123, -47, -117, 23, 15, -107, 76, -44, 9, 38, 104, -107, -1, 59, 79, 93, -23, 63, -116, -126, -35, 120, -120, -48, 97, 121, 102, -34, -105, -36, -35, -100, 45, -24, 51, -67, -3, 0, 17, -121, -90, -6, -100, 37, -75, 107, 2, 30, 43, 15, 32, -120, 7, 40, -40, -24, 33, -66, 70, 56, 26, -93, 84, -56, 12, 7, 5, -119, -121, -106, -112, -82, 16, -83, 83, 69, -104, -42, -29, 67, 101, -125, 75, -20, 43, -92, 84, -52, -30, 26, -124, 125, 61, 88, -59, -55, -32, 74, -45, -25, 96, -29, 21, -15, 16, -23, -74, 41, 63, 26, -20, 36, 29, -72, -112, -55, -36, 100, 21, 62, -2, 26, 59, -69, -14, -128, 5, 82, 74, 88, -70, 43, -69, 79, -100, 76, -72, -46, -11, 119, 108, 97, 27, 10, -103, 43, 83, -11, 15, -24, -76, -115, -126, 111, -55, -11, 112, 78, -57, 58, 38, 1, -27, 97, -47, 1, 45, 9, 84, -94, 1, 64, -124, -100, -54, -99, 72, -99, 19, -41, 6, 71, -27, 8, 54, 46, 125, 38, -4, -59, -31, -94, 70, 70, -125, -105, -56, 49, 33, -100, 83, -94, 92, 87, -66, -89, 117, -122, -60, 8, -34, 74, -49, 67, -45, -123, -15, -48, 44, 109, 21, -115, -113, -36, 83, -110, -13, -101, 67, -108, -73, 23, -74, -108, -18, -11, -69, -29, -5, -1, 107, 89, -54, -70, 28, 29, -64, -115, 109, 108, 122, 3, 121, -119, 95, 76, -100, -46, 104, 95, -25, -97, -10, 29, -77, 101, -110, -18, -56, 14, 110, -76, -25, -72, -18, -124, 85, 46, -111, 66, 26, -116, -59, 19, -107, -92, -32, -79, -9, -56, -111, 94, -25, 7, -5, 27, -20, 14, -119, 53, -100, 119, 105, 3, -81, -41, 7, -124, -122, 25, 71, 32, 37, -116, -76, 58, -79, 20, 108, 40, 92, 125, 6, -61, 4, -127, 94, 113, 15, 104, 38, 43, 95, 15, -81, -113, 102, 54, -109, 108, -49, 90, 13, 116, 103, 65, 47, -104, -43, 27, 64, -79, 24, -58, -12, -100, -57, -45, -115, 87, -69, 51, 2, -102, -62, 49, -87, -87, -24, -67, -107, 55, -105, 34, 44, 126, -29, -37, -106, 56, 118, 86, 105, 14, -100, -34, 42, -28, 49, 56, -69, 108, -21, 61, -122, 46, -17, -80, 87, 87, -19, 108, 14, 4, 15, -70, 3, 114, 21, 25, 43, 11, -16, 20, -103, 12, 114, 68, 112, 35, -4, -85, 15, 103, 105, 22, 21, -40, 70, -20, -81, -77, -39, 61, 55, 104, 120, -70, 90, 13, 84, 5, -103, -60, -102, -78, 80, -116, 118, 65, 48, -14, 108, -65, -38, 85, 85, 111, -83, 27, -36, -36, 78, 53, -102, 6, 29, -110, 64, -9, 31, 20, 125, 56, 88, -105, 107, 41, -93, 97, -22, 83, -44, -42, -109, 46, -84, 104, 29, -39, 4, 121, 54, -46, 46, 80, 88, -53, 98, 25, 67, 1, -83, 64, -70, -122, 87, -91, 47, 122, -122, -103, 78, -38, -17, 97, -120, 27, 73, 38, 117, -51, 31, 43, 32, -50, -5, -8, 25, -35, -111, -36, 94, -65, -100, -104, -59, 115, -67, 116, 110, -60, -115, 60, 30, -4, 29, 39, -104, -26, -51, -115, 52, 108, 56, -44, -70, -77, 76, 84, 16, 94, -80, -18, -99, -51, 7, -30, -64, 68, -42, -82, -120, -29, 106, 39, 95, 7, -50, 119, 110, 27, -124, 34, 7, 60, 118, 66, 111, 66, 22, -1, 32, 70, 110, 61, -109, -11, -97, -44, -71, -11, 2, -62, 88, -19, 105, 56, 116, -73, 47, 98, 82, 52, 4, -39, -16, -6, -101, -32, -67, 49, 95, 93, -8, 77, 27, 11, -62, 58, 95, -4, -80, -30, 62, -120, 79, 39, 64, 67, 94, -16, 38, 48, -92, -86, -119, 20, 37, -91, 116, 98, 86, 84, 63, -50, 33, -38, 90, 100, -107, 57, -32, -59, -101, -98, -51, 106, 69, -114, 46, 35, -2, -44, -45, 34, -2, -36, -74, -93, 1, -85, -123, -40, 127, 69, 38, 32, -97, 0, 4, -76, -70, 100, -7, -43, -126, 71, -64, 71, 85, 110, -22, -45, -62, 61, 117, 64, -102, -85, 100, 27, -42, 105, 115, -43, 46, 26, 118, 78, -102, -6, -126, -44, -33, -4, 42, -31, -61, 106, -87, -104, 88, 19, -21, -102, -47, -32, 90, -21, 11, 62, -122, 98, 40, 122, -73, -42, 20, -83, -92, 46, 40, -89, -125, -121, 35, 45, -24, 102, 23, 17, 126, -17, -91, -23, 9, -10, 73, -29, 97, -44, -94, 103, -74, 74, 97, -18, -96, -11, 27, -59, -92, -61, -20, -89, -54, -113, 84, 51, 117, -21, -60, 115, 90, -23, -36, -29, 95, -91, 70, 64, -7, 104, 40, 48, 50, 9, -98, 83, 127, 57, -104, -93, 125, 4, -54, -57, 19, -98, 122, 8, 9, -65, -5, -29, 40, 87, 70, 8, 124, 12, -56, -11, -11, 112, -91, -89, -6, -61, 122, -7, 125, -110, 28, 122, 22, 102, -63, -87, -124, -68, 49, 13, -5, -84, 112, -93, -125, 54, 43, 127, -62, 116, -11, 55, 100, 26, 95, -34, 94, 89, 87, 91, 108, -13, 85, 2, -39, -106, 44, -35, -46, -35, 106, 77, 10, 90, 113, 13, 16, 28, 13, 83, 16, -126, 10, -11, 28, -23, 83, -6, -61, 43, -43, -81, -98, -86, 49, -8, -63, -35, 85, 19, 59, 64, -31, -59, 26, -46, 82, -85, 110, -33, 126, -1, -31, 8, 116, 126, 114, 71, -8, -75, -14, 78, -28, 17, 120, -107, -119, -71, -13, 94, 77, -82, 30, -82, -13, -71, 0, -59, -28, -18, 37, -30, 109, -122, 106, 97, -124, 92, 41, -3, -111, -101, -53, -11, 44, -61, 11, 53, -3, 126, 20, -54, -84, -78, -8, 31, -21, 120, 100, 79, -26, 9, -79, -44, 16, -100, -75, 20, 120, 94, -111, -118, 122, -36, -1, 38, 32, -118, -36, -99, -120, 112, -25, -76, -94, 95, 83, 14, 87, 56, -35, -67, -63, 15, 17, 81, 43, 71, -26, 35, 37, -9, 45, 31, 84, -83, -58, -12, -73, 34, 17, -64, 18, 120, -12, 52, 87, -56, -62, 46, -128, 32, 107, -63, -81, -3, -109, 90, -60, -7, -3, 105, 112, -85, 9, 68, -40, 79, -72, 15, -15, 73, 79, -125, 65, -60, 55, 24, 12, 122, -58, 12, 26, -78, 77, 73, 47, 96, 35, 115, -39, -96, 92, -54, -53, -27, -114, 35, -76, -57, -77, 37, -112, -126, 40, 82, -58, -32, -22, 82, -38, 49, -34, 116, 99, -84, 61, 18, -116, -32, 5, -26, 0, -31, 48, 76, 71, 62, -17, 123, -123, 34, 33, -106, 37, -55, 104, 107, 41, -46, 62, -125, -125, -100, 119, 102, -56, 52, -8, -43, -108, 125, 59, 21, -33, -21, -31, -90, -87, 80, -95, -81, -13, 66, -59, -104, -116, -83, -125, 53, -1, 65, 57, 3, 94, 48, -23, -90, -27, 98, -5, -7, 95, -74, -114, -66, 33, -17, -28, 75, -64, 6, 122, 51, -56, -65, 75, -44, -20, 78, -118, 107, 16, 67, -18, -18, -13, 88, 20, 88, 58, -112, -46, 25, -58, -32, 88, 104, 80, -68, 51, -112, 66, 45, 67, -117, 108, 14, -33, -40, -36, -23, -61, 108, -84, 50, -38, 32, 10, 111, -8, -60, 127, 74, 93, -59, -85, 53, -83, 123, 114, 96, -117, 52, 13, 78, 63, -7, -36, -97, 81, 56, 8, -107, 37, 53, 71, 127, -43, -47, 110, 77, 21, 109, 24, -14, -77, 67, -88, -32, 62, -102, -63, 73, 78, 78, 23, 14, -56, 115, 45, -103, 43, -75, -82, -48, 106, 117, -48, -65, -58, -66, -115, 91, -84, 37, -50, -33, -24, -10, 63, -90, 16, -128, 111, -34, 79, 6, 108, -105, -7, 25, -80, -92, 79, -33, -11, 57, -44, 69, 121, 27, -125, -122, -10, -81, 43, 68, 14, -109, -70, -50, -71, 74, -50, -88, -87, -99, 46, -107, -76, -89, 47, -27, -53, -2, 68, 64, -73, -104, 5, -80, 51, 9, -74, -86, 56, 97, 110, -57, 116, -87, 21, -83, 115, 99, -43, -100, -127, -125, -78, -75, -86, 97, 26, -10, -33, -34, -74, 22, -9, 60, 71, -86, -59, 125, -44, 125, 95, -61, -60, 83, -20, 89, -127, -33, 61, -42, -4, 62, -38, 46, 115, 4, 15, 14, 122, 110, 108, -79, 4, -29, 109, -53, 14, -78, -55, 98, -81, -88, -91, -12, 123, 17, -51, 124, 113, -118, -45, -19, 72, 45, -101, 60, -79, 42, -54, -84, 24, -74, -35, -100, 26, -54, -24, -88, -4, 49, -118, 43, 89, -80, -97, 84, 65, -19, 81, 50, -9, -92, -97, -64, 81, -70, 124, -126, 100, -58, -82

);
    signal scenario_output : scenario_type :=(6, 12, -2, 58, 90, -97, 1, 45, -100, 23, -52, -68, -21, 59, 127, -44, 2, -70, -33, -18, 60, -6, -128, 127, 12, -79, 44, 63, -12, -112, 122, 100, -128, -55, 44, -6, 43, 13, -96, -2, 49, 27, 42, -23, 78, -2, -16, 50, -42, -81, 63, -11, -79, 87, -73, -12, -23, 2, 16, -27, 47, -57, -43, -47, 60, 117, -86, -71, -3, 15, 37, -5, 33, -117, 21, 81, -90, -6, -1, -79, -58, 70, 86, -2, -38, -103, 12, 112, 33, -128, -29, 116, -26, -127, 97, 24, -128, 42, 127, -12, -128, 53, 10, 71, 71, -128, 38, 13, 23, -12, -32, -44, -76, 81, 127, -2, -52, -32, -5, 12, -1, -68, -6, 2, 2, 37, 37, -5, 48, -28, 11, 45, -6, -128, 2, 97, -123, 11, -22, -45, 7, 121, 23, -101, 24, 17, 93, 90, -44, -91, -11, -15, 16, 97, -64, 10, -42, -128, 55, 16, 27, 36, -70, 50, 59, 66, -69, -8, 47, -81, 79, 23, -128, -31, 121, 1, -43, 34, -23, -57, 123, 78, -106, -34, 60, -118, 3, 28, -80, 127, -3, -64, 15, -23, -42, 108, 11, -80, 65, 69, -6, -52, -39, 52, 50, -119, -59, 37, 95, 29, -49, 39, -24, 63, -26, -121, 127, 92, -128, 50, 70, -96, -22, -68, 76, 48, 7, -109, 21, 42, -6, -15, 18, -58, -100, 103, 0, -44, 91, 63, -23, -128, -11, -16, 102, 74, -128, 68, 32, -95, 90, -50, 28, 13, -90, 75, 95, -113, 0, 86, -37, -16, -68, 12, 100, -31, -101, 127, 57, -42, 15, -78, -128, 13, 101, -75, 101, 66, -38, -64, 23, 17, -85, 22, 42, -15, -98, 1, 91, -128, -48, 81, 27, -1, 65, -70, -2, 122, -128, -58, 127, -112, 37, 119, -128, -58, 95, -37, -128, 86, 97, -128, -31, 43, 87, -39, 57, -43, -6, 117, -128, -66, 43, 85, 66, -111, 64, 52, -128, 127, 109, -44, -128, 32, 106, -95, -55, 42, 65, -48, -69, 26, 13, 12, 37, -96, 24, 65, -108, 6, 26, -50, 53, 16, 21, -76, -38, 54, -12, -28, -16, -17, -43, 15, -16, -73, -45, 103, 106, -128, -59, 66, 24, 91, -118, -49, 24, 106, -34, -49, 79, 0, 53, -63, -96, 107, 55, -128, 26, 74, 0, -22, -78, 8, 3, 79, 50, -73, 5, 21, -32, -87, -45, 44, 13, 11, 109, 8, -80, 103, 96, -31, -71, 12, 102, -32, -76, 23, 17, -80, -34, 49, 71, 0, 8, 65, -97, -52, 23, 107, -85, 21, -10, -100, 33, 12, 47, 92, -6, -43, -1, 119, 59, -106, -44, 47, -87, -91, 85, 109, -57, -3, 127, 3, -128, 22, 102, -80, -60, -8, 54, 31, 127, -6, -79, -34, 37, 103, 3, 0, 28, -7, -58, -24, -60, -71, 32, 28, -47, 86, -58, -53, 70, -65, -17, 65, 70, 29, -24, -128, 73, -1, -127, 127, 1, -68, 80, 28, -128, -28, 80, -80, -6, 52, -74, -58, 127, 73, -59, -66, 23, 78, 12, -123, 64, -36, -26, 127, -128, -21, 127, -121, 6, 0, -87, 38, 109, 127, -128, 17, 68, -36, -71, -73, 47, 29, 2, -12, 127, 78, -113, -16, 42, -68, 55, 54, -73, 18, 24, -15, 127, -57, -86, 112, -45, -34, 100, 50, -106, 2, 59, -128, -1, 127, -128, 12, -1, -96, 127, -86, 33, 11, -71, 45, -23, -45, 113, 36, -57, -59, 73, 44, -87, -22, 0, 65, 76, -98, 1, 2, 102, 10, -128, 90, 18, -48, 50, 27, 10, -11, -3, 12, 29, -109, 70, 127, -128, 5, 43, -47, 79, -80, -117, 24, 73, -1, 57, -47, -47, 29, -11, 23, 50, 5, -106, 103, 92, -86, -44, -32, 100, 64, -48, -66, 7, 10, -59, -128, 48, -6, 23, 75, -76, 43, 70, -128, -71, 127, -50, 13, -28, -11, 6, 32, 127, -128, -39, 86, -16, 27, 21, -95, -21, 23, -128, 15, 45, -12, 24, -103, -128, 102, -16, -12, 95, 63, -59, -8, 24, -58, -24, 27, -103, 11, 49, -111, -64, 17, 127, 52, -128, 59, 10, -128, 95, 57, 11, -55, -70, 68, 15, -69, -47, 50, -96, -90, 127, 42, -128, 34, 13, 42, 11, -55, 44, -95, 29, 95, -107, 6, 11, -36, 13, 33, -21, -90, -22, 39, -116, -60, 121, 76, 2, -124, -5, 107, -78, -57, 11, 8, -73, 58, 21, -29, -7, -91, 95, -7, -128, 39, 8, 78, -48, 54, 80, -38, -43, -75, 32, 17, -2, -43, -16, 31, 28, -54, 1, -17, 86, -34, 23, -18, 53, 12, -18, 13, -44, 43, 15, -18, -114, -90, 90, 13, 101, -27, -128, 90, 71, 28, -91, -44, 15, 69, 101, -5, 2, -95, 27, 55, -98, 18, 68, -75, 64, 16, -29, 7, -73, 36, -1, -8, 63, 33, -5, -32, 36, 10, -128, -2, 71, -54, 65, 36, 2, -8, -85, 36, 71, 58, 43, -36, -98, -23, 106, -86, 23, 43, -45, -58, -74, 127, 44, -43, 6, -74, -24, 54, 113, -53, 21, -12, -57, 54, 32, 80, -5, -59, -57, -48, 49, -3, 93, 66, -58, 0, 31, -44, -93, 16, 71, -32, -28, -17, 121, 92, -128, 85, -49, 16, 0, 2, -26, -26, 26, 37, 22, 50, -52, -23, 127, -54, -38, 54, -103, -47, 64, 107, 21, -58, -52, -39, 106, 31, -91, 48, -10, -17, 80, -28, -31, 91, 109, -91, -128, 127, 85, -128, 21, 60, -8, -36, -108, 1, 27, -33, 69, 60, -103, -22, 32, 18, 50, 87, 21, -49, -63, 39, 66, -32, 1, -128, -57, 127, -53, -54, 92, 59, -42, -86, 7, 0, -112, 100, -49, -52, 33, 50, -21, -58, 127, -39, -48, 16, 98, -58, 0, 2, 12, 55, -128, 45, 92, -87, -8, -76, -91, 113, -5, 65, -23, 33, 33, -103, 102, -5, -21, 86, 13, -52, -128, 43, 106, -64, -128, 66, 95, -128, -64, 127, 65, -93, -11, 42, -128, -10, 127, -103, 49, 107, -48, -128, 24, 16, -57, 75, 21, 78, -34, -76, 55, 10, -65, 26, -21, -3, 60, -85, 24, 114, 23, -87, -93, 63, -32, -23, 0, 121, 28, -128, 112, 11, -101, 86, 38, -22, 111, 50, -121, -38, 3, 113, 86, -93, -36, -71, 122, -26, -124, 116, 118, -128, 59, -6, -36, -2, -18, 98, 65, -21, -58, -21, 21, -2, -128, -74, 127, 92, -54, -127, -85, 127, -64, 31, 43, -92, 117, -53, -65, -38, 93, 21, -128, 123, 24, -43, 68, -3, -123, 17, 24, -128, 28, 55, 23, 8, -48, 17, -11, -73, 70, 37, -123, 57, 38, -48, -43, 0, 96, 5, -71, 11, -109, 3, 85, -50, -49, 15, -23, 24, 3, -128, -73, 43, 100, 65, 22, -128, -29, 39, -1, 7, -75, 93, 13, -5, 12, 1, -15, -24, 37, 111, -64, -38, 102, -117, -37, 63, 76, 71, -109, -32, -31, -3, 124, 34, -117, 12, 108, -10, -128, -8, 28, -22, 29, 53, 108, -6, 23, 59, -42, -116, 33, 91, -17, -80, 24, -90, 12, 71, 13, -107, -117, 127, 2, -22, 17, -59, -21, -8, -38, 11, 95, -63, -39, 95, -18, -111, -26, 54, -38, 108, 54, -34, 18, -78, -65, 55, 29, -81, -6, 75, -11, 10, 37, 42, -22, -76, 12, 127, 26, -57, -29, -12, 75, 64, -117, -58, -13, 33, 111, -86, -34, 28, 97, -66, -16, 0, 18, -17, -50, -16, 68, 70, -37, -70, -21, 127, -33, -38, 74, 24, 37, 11, -128, 0, 108, -85, -91, -42, 1, 29, 48, 79, 27, -49, 65, -21, -17, 53, -28, 65, 5, -128, 21, -1, -31, 116, 86, -75, -102, 44, 0, -31, 66, 32, -64, 17, 127, -39, -74, 118, -42, -34, 0, 16, 69, -128, -118, 81, 98, -11, -49, -31, 47, 87, -86, 3, 23, -116, -38, 101, 44, -69, -109, -23, 127, -57, -34, 111, -45, -122, 71, 109, -21, -127, 11, 78, -80, 28, -34, -97, 47, 91, 5, -103, 42, 127, -128, -68, 54, 28, 0, -54, 127, 6, -112, 119, -18, 8, 11, -13, -123, -52, 127, 31, -42, -58, -2, -71, -17, 127, -54, -1, 29, -16, 50, -127, -12, 121, -78, 10, -48, -26, -54, -26, 10, 31, 39, 22, 8, 81, -22, -80, 18, -31, 1, -10, 86, 114, -116, -112, 117, 26, 21, -50, -106, 103, 21, -128, 90, -3, -108, 49, 127, -47, -28, 127, -47, 0, -48, 13, 52, -39, -76, -60, -39, 102, 39, 11, 16, -21, -109, -1, 36, 90, 60, -100, 15, -50, -31, 52, -45, -2, 70, -100, 1, 31, -108, 5, 43, 39, -10, -37, 29, 90, 12, -42, -6, 108, -59, 42, 52, -128, 7, 121, -58, -64, 52, 127, -1, -8, -11, 2, -22, -75, -43, -10, 127, -36, -36, -21, 33, 88, -92, -112, 39, 121, -37, 2, 28, -45, 12, 93, -49, -7, 15, -76, 60, 36, -122, -54, 58, 65, -85, -100, 21, 49, 24, -64, 65, -42, -53, 90, -112, 52, 93, -101, -24, 107, -108, -128, 92, 81, 74, 10, -102, -22, -15, -8, 24, 39, 70, -114, -8, 17, -13, -38, 101, -21, -73, 127, -32, -128, 69, 53, 48, -55, 5, 11, -107, 96, -3, -45, 1, -43, -2, 76, 47, -50, -109, -39, 39, -26, 42, -18, 23, -2, -28, 95, -13, 53, 10, -13, 50, 48, -128, -12, 22, 65, -52, -50, 127, -26, -108, -22, 127, 23, -128, 59, 3, -54, -32, 55, 53, -42, 26, -121, 5, -32, 3, -38, 50, -15, -23, 93, -124, 55, 26, -69, 91, -15, 34, 2, 8, -103, 10, 107, -48, -128, 31, -11, 0, -31, -92, 106, -42, -53, 127, 76, -119, -31, 91, -98, -15, 34, 5, 13, -107, -81, -1, -3, 100, -16, 28, 76, -91, 28, 48, -108, 85, 27, -90, 53, 5, -23, -58, 13, -90, -32, 124, -10, -97, 58, 90, 22, -106, -18, 69, -32, 11, 15, -49, -64, -117, 31, 23, -8, 7, 85, 38, -106, -2, 2, -17, 12, 127, 34, -22, 34, -7, -75, -91, -50, 12, 8, 127, 23, -42, 38, -124, 22, 66, 23, -95, -17, 24, -37, -59, 65, 12, -8, 97, -42, -37, 45, -37, -57, -32, -8, 7, -8, -74, 96, 50, -114, 95, 1, -36, 42, -116, 55, 12, -16, 48, -48, -47, -60, -55, 92, -48, -11, 49, 78, -63, -122, 127, 74, -44, -74, -48, -5, 93, 10, -109, 8, 117, -65, 42, 47, -11, 81, -95, -114, 118, -33, 34, 17, -64, -29, -45, 85, 71, -26, -33, 39, 7, -75, 0, -5, 26, 65, -43, -55, -57, 44, 65, 5, -31, -68, -59, 6, 23, 22, 28, -75, 38, 32, -26, -54, 12, 60, -1, -91, -78, 15, -17, -59, 118, 97, -98, -29, 48, -91, -78, 127, 69, -43, -2, -75, -59, -52, 108, 78, -60, -38, -112, 29, 3, 58, -55, -117, 127, 119, -71, -122, 0, 108, -47, -79, 69, 52, 23, -101, 13, -64, -69, 116, 91, -103, -96, 59, 39, -17, 3, 10, 118, 6, 10, -53, -68, 127, -34, -114, 127, 91, -101, -60, 60, 49, -6, -66, -10, 48, 28, -48, -5, 97, 34, -93, -122, -27, 127, 33, -100, 119, 13, 6, -49, -111, 127, 15, -128, -21, 101, 95, 15, -8, -128, -34, 70, 26, 11, 28, -102, -73, 10, 91, -7, -88, 27, 47, 0, 122, 50, -112, 42, 118, -128, 22, -1, -118, 69, 17, -3, -27, 0, 43, 127, -29, -22, 11, 47, -21, -95, -22, 80, 31, 15, 42, -87, 33, -108, -34, 124, -45, 8, -29, -43, -71, 1, 127, -75, 39, -48, -48, 127, -101, -13, 90, -78, -49, -32, 0, 106, -11, -52, 7, -95, 13, 60, 15, -1, -12, -28, -12, -7, -8, 127, 60, -113, -42, 57, 29, -53, 39, -28, -60, 127, -75, -108, 111, 50, -26, 79, -21, -128, 58, 127, -113, -124, 92, 102, -11, 45, -128, 24, 6, -106, 127, 79, -59, -114, 22, 0, 29, 10, -16, 124, -48, -63, 127, 8, -21, -50, -23, -11, -6, 2, -2, 76, -5, 57, -17, 32, 73, -114, 26, 91, -60, -43, 33, 74, -42, 3, 43, -22, -128, -90, 127, -31, -13, 64, 29, -68, 43, -24, -49, 3, -10, 81, 29, -27, -57, 64, -26, 24, 86, -28, -59, -92, -21, 2, -6, 127, -22, -98, 127, -6, -50, 54, -6, 68, 90, -128, -116, 127, -1, -28, -48, 38, 22, 12, -18, -2, 45, -13, 10, -2, -12, 127, 17, -87, 100, 0, -128, -57, 101, 127, -96, -128, 47, 95, 75, -81, -6, -48, -53, 21, 100, 11, 7, 91, -5, -22, -91, -73, -6, 98, 36, -50, 27, 88, 17, -70, -45, 86, 5, -128, 76, 109, -128, -73, 90, -27, 42, 28, -66, 124, 0, 0, 106, -2, -86, -12, 6, 1, 26, -29, -76, -70, 117, 64, -13, -43, -121, -8, 52, 60, -16, -66, 34, 43, -26, 71, -15, 3, -96, -29, 98, -64, -38, 45, 127, 8, -128, 21, 42, 59, -59, -3, -21, -79, 92, 127, -8, -59, -45, -70, 32, 113, -23, 36, -42, 1, 78, -26, -23, 12, -68, -81, 127, 5, -66, 101, -119, -12, 70, -45, 13, 39, -79, 3, 96, -18, -32, -27, -48, 97, 15, -47, 10, 44, -39, 0, 15, 68, -57, 22, 52, -95, -69, 43, 109, 0, -74, 42, -44, 26, -34, 1, 36, -86, -3, -22, 93, 75, -79, -128, 37, 127, -45, -128, 43, 112, -31, 27, -16, -36, 39, -101, -101, 127, 54, -22, -28, -128, 49, 124, -128, 44, 95, -91, -49, -65, 106, 10, -124, 54, 54, 49, -28, 38, 37, -16, -26, -109, 63, -33, 52, 52, -103, -58, 44, 127, 31, -13, -128, -31, 127, -122, -17, 79, -13, 44, -15, -87, -78, 55, 85, -54, -69, -59, 34, -18, 100, 124, -128, -13, -23, -54, 48, 49, 0, 60, 22, -81, 78, 37, 17, 1, -29, -8, -53, 5, 47, 107, 33, -63, -12, 2, -65, -71, 121, 86, -127, 42, 74, -66, -23, 59, 11, -27, 78, 1, -128, -33, 117, 50, -26, -39, -60, -24, 127, -1, -50, -2, -7, 13, 111, 92, -32, 11, 7, -91, -36, 80, 65, 5, -128, -73, 98, 27, 33, -18, -107, 91, 59, -18, -33, -80, -28, 79, 6, 44, 47, -74, 8, 6, -70, -55, -13, -52, -11, 2, 32, 87, -113, -13, 124, -98, 47, 3, -17, 49, -5, 32, -57, -59, 43, 85, -26, -16, -32, 32, 16, -121, 8, 57, -81, -29, 11, 79, 31, -29, -95, -49, 87, -29, 70, -6, -75, 87, 6, 60, -81, 53, 63, -109, -16, -27, 6, 127, 68, -55, -10, -28, -128, 29, 37, -31, 116, 18, -128, 32, 17, -45, 98, 54, -87, -28, 78, -5, -128, -28, 87, -24, -6, -5, 64, 91, -87, 60, 24, 33, -5, -121, 34, 44, 24, 22, 1, -36, -93, 93, -54, -42, 13, 73, -16, -38, 33, -74, -13, 70, 8, 18, 13, -28, 3, -98, -74, 127, -90, -16, 127, -86, 17, -43, 11, 32, -128, 66, 6, -49, 108, -36, 43, 91, -128, -91, 80, 70, -29, -128, 26, 8, 87, -10, 11, 58, -76, -73, 38, 31, 44, -38, 0, 31, -50, 0, -91, 10, 13, -52, -49, -33, 127, -37, -78, 17, 48, 118, 36, -11, -22, -113, -118, 96, 53, 28, -42, -128, 7, 7, 92, 0, 0, 58, 63, -60, -74, 23, -39, 118, 87, -123, -93, 79, 36, -55, 47, 74, -116, -28, 114, -107, -128, 127, 106, -111, 24, -71, -28, -17, -32, 31, -6, 102, 59, -121, -74, 15, 79, 17, -63, 31, 95, -18, -86, -3, 122, 97, -128, 58, 33, -2, -76, -66, 127, 57, -128, 27, 15, -16, -43, 13, -15, -18, 86, 53, -3, -21, -107, -37, 28, 7, 109, 70, -42, -7, 55, -98, -48, 127, -69, -128, 127, 28, -79, 96, -47, -47, 70, 0, -96, 58, -16, -80, 7, 100, -57, 33, 45, -128, -33, 87, 10, 39, -38, 18, 21, -119, -24, 3, 17, 80, -7, -43, 127, 47, 17, -81, -114, 122, 93, -74, -15, -58, 42, 127, -128, -128, 127, 65, -128, -39, 16, 101, -50, 7, 91, -17, 24, 12, -44, 33, -102, -22, 127, 8, -128, 29, -42, -68, 100, 63, 11, -114, -112, 108, 22, -92, 113, -2, 5, 119, -96, 11, 23, -95, 8, -42, 106, -15, 2, 48, -128, 121, -3, -128, 127, 18, -2, 68, -58, -79, 15, -13, -17, 39, -107, -128, 127, 121, -128, -23, 107, -42, -43, -26, 60, 80, -101, -10, -49, -43, 48, 7, 24, 54, -2, 127, 64, -128, 88, 34, -66, 73, -114, -32, 124, -43, -28, 73, -55, 23, -2, 58, 117, -76, -128, 63, 32, -47, 0, -5, 43, -1, -27, 36, 21, -42, -3, -48, -7, 29, 17, -86, -50, 102, 15, -127, -54, 17, 124, 2, -8, 112, -116, -6, 63, -63, 3, 108, 23, -24, -74, -45, 2, 95, -39, -111, 85, 127, -23, -122, 48, 24, -29, 127, -69, -128, 36, 52, 5, 111, 23, -13, 22, -38, -50, 97, 31, -78, 26, -57, -52, -36, 71, 65, 5, 0, -54, -87, 16, -47, -10, 12, -10, 116, -73, -28, -43, -24, 127, -69, -93, 47, 114, 43, -23, -116, 26, 38, 2, 1, 11, -79, -2, 53, 16, -7, -79, 13, -64, -50, 127, 38, -68, -44, 17, 76, -127, 6, 21, 43, 73, -103, -86, 71, -27, 68, 70, -31, -68, -38, 22, -45, 78, -32, 38, 64, -10, -50, -75, 123, 32, -128, 26, 127, -38, -128, 107, 32, -7, -70, -36, 96, 1, 12, -50, 26, 49, 50, -34, 11, -18, -2, 102, 6, -47, -33, -42, -26, 92, 13, -102, -10, 81, 59, -65, 73, 44, 7, -69, -100, 127, 7, -33, -39, -114, 112, 101, -95, -33, 96, 52, -86, -86, 39, -26, -101, 15, 109, -12, 75, -73, -64, 33, 17, 127, -63, -85, 60, -22, 23, 98, -88, -81, 95, 48, -60, 8, 12, 39, 111, -88, -18, 54, 23, -29, 38, 58, -45, -48, 97, 0, -92, 1, 44, 81, -86, 33, -31, -11, 127, -38, -92, -75, 75, 119, -79, 2, -69, -12, 12, 50, 32, -36, -69, -78, 127, 86, -49, -95, -78, 76, 81, -55, 48, -49, -88, -5, 127, -5, -49, 111, 6, -128, 65, 50, -22, -23, -79, -39, -27, 112, 124, -26, -102, -79, 114, -3, -128, 95, 78, -74, -24, 24, 66, 127, -75, -31, -45, -49, 127, 38, -128, 32, 86, -103, -49, 95, 47, -15, 1, 8, -80, 11, 12, -5, 66, -91, 18, 71, -26, -98, 28, 85, -103, -80, 86, 37, -128, 70, -43, 26, 78, -128, 48, 7, -54, 113, 50, -16, -79, -60, 22, 34, -101, 68, 0, -1, -31, -116, 122, -48, -15, 98, 45, 33, -128, 15, 106, -128, 34, 93, -128, -39, 127, 31, -63, -92, 28, 39, -78, -39, 127, 58, -34, -122, 12, 13, -114, 127, 12, -23, -88, 48, 43, -10, 52, -106, -3, 1, -33, 0, -59, 31, 95, -118, -49, 60, -10, -52, -53, 109, 39, -96, 53, 36, -18, 13, 60, 22, -45, 127, -31, -102, 127, 42, -124, 63, -31, 69, 12, -34, 37, -15, -12, -23, 63, 70, -128, -60, 48, -36, 127, 37, -128, 15, 107, -26, 0, -29, 26, 91, 44, -34, -22, 12, -128, 70, 24, -128, 111, 48, -7, -49, -81, 8, 102, 117, -128, -5, 22, -78, 113, -33, -8, 106, -48, -80, -55, 127, 1, -60, 63, -66, -45, 49, 123, -38, -74, 11, 27, 127, 28, -128, -37, 127, -32, 32, 63, -119, -2, 97, -42, -90, -50, 0, 27, 76, 31, -60, 28, 65, 32, -128, 29, 123, -108, -22, -52, 13, 103, -54, -12, -1, -13, 85, -75, 3, 87, -1, 42, -116, -18, 29, -26, 43, -21, -8, -55, -103, -17, -16, 127, 127, -128, -7, 117, -64, -81, 96, -59, -116, 70, 103, -2, 24, -8, -26, -1, 108, -38, -96, 22, 118, 48, -34, -13, -88, 6, -60, 6, -64, -48, 116, 75, -68, -92, 57, 65, -37, -65, 36, -17, -26, -36, -128, 28, 127, -47, -2, 37, -33, -111, -73, 116, 127, -128, -34, 80, 43, 36, -128, 29, -22, -128, 127, 87, -107, -2, 36, -93, -36, 86, 87, -95, -109, 127, 48, -8, -74, -69, 79, -98, 0, 122, -13, -60, 31, -59, -116, 127, -13, -45, 108, -26, -39, 47, -75, 70, -5, -6, -52, -11, 66, -122, 91, 73, -3, -36, -50, -26, -74, 39, 50, 58, -36, -76, 49, 5, 36, 49, 81, -7, -7, -7, 16, -59, -96, -5, 21, 96, -64, 0, 52, 12, 32, -54, -27, 59, 85, 34, -16, 0, -101, -80, 88, 39, -43, 87, 13, -15, -42, -15, 6, 127, 91, -6, -111, -121, 17, 90, 91, -76, -88, 6, 127, 58, -100, 74, 90, -24, -65, -43, 2, 10, 10, -127, 81, 102, -70, -79, -49, 86, 17, -73, 34, -6, -48, 106, -11, -60, 15, -55, 58, 42, -80, -3, 127, -23, -128, 108, -17, 3, 11, 15, -15, 32, 45, -128, 21, 6, -12, -59, -43, 34, 43, 108, -22, -15, 11, 16, -90, -107, -6, 127, 49, -119, -33, 48, 53, -26, -60, 88, -52, -17, 71, -36, 3, -36, 48, -26, 0, 2, -54, -74, 49, 123, 0, -128, -7, 65, -100, -87, 127, 27, -128, 52, 107, -33, -97, 24, 127, -22, -86, -29, -8, 127, 45, -36, -49, -18, -11, -17, -3, 111, 21, 13, 54, -92, -81, 57, 127, -68, -58, 91, -7, -37, -54, -36, 124, -36, -43, 63, -27, 6, -18, -48, -6, -90, -32, -45, 69, 69, -117, 53, -17, -43, 57, -119, 60, 91, -92, 34, -92, -98, 127, 76, -22, 50, -128, -11, 44, 16, 18, -119, 74, 8, 29, 15, -47, -33, 1, 10, -101, -63, 75, 57, 27, -86, -7, 58, 36, -112, -60, 127, -73, -123, 87, 123, -124, -17, 79, -48, -11, -55, 50, 11, -13, 50, 59, -73, -119, 116, -50, -42, 127, -6, -128, 57, 107, -33, -80, 7, 73, -128, 16, 31, -98, 73, 0, -3, 1, 90, 81, -60, 22, -63, 1, -3, -128, 95, 100, -128, -10, 79, -15, -43, -63, 38, -15, -92, 36, 101, -114, -44, 127, -128, 16, 13, -44, -12, 21, 93, 44, -73, -85, 97, 59, -113, -60, 127, -49, -98, 31, 127, -69, 45, 63, -102, 75, -109, 24, 60, 22, -100, -119, 127, -49, -128, 58, 102, -31, 49, -2, 43, 112, -117, -34, 36, -10, -128, 11, 127, -113, 12, 76, -128, 48, -15, -11, 71, -95, 1, -1, -38, 78, 13, -57, 59, 16, -28, -33, 37, -11, -5, 71, -55, 95, -13, 10, 52, -114, 12, 33, -6, -3, -45, 80, -7, -29, 37, 74, 10, 7, -124, 22, 55, -78, -44, -38, 127, 38, -107, -21, 58, 22, -1, -7, -58, -128, 54, 3, -48, 15, 48, 79, -38, -6, -34, 3, -68, 31, 47, -26, 8, -44, -12, -69, -69, -47, 90, 15, 22, -47, 23, 49, 6, 11, -93, -21, 76, -91, 12, -1, -42, 52, -57, -28, 55, 85, 90, -43, -59, 22, -17, -17, 8, -21, 88, 53, -101, -18, 122, -111, -34, 117, -28, -39, -6, -69, -29, 79, 16, 98, 24, -34, -45, 0, 69, -21, -95, 23, 127, -17, -128, 0, -6, 34, 92, 49, -108, 42, 18, -128, 127, 98, -55, -75, -57, -32, 31, 27, -3, 37, -50, -93, 33, 78, 42, -93, -76, 127, 65, -128, -7, 113, -28, -47, -27, -50, 33, 63, -59, 64, 76, -128, 47, 52, -6, -60, 49, -6, -2, 34, -103, -23, 119, 44, 23, -36, -15, 103, -90, -65, -7, 101, -3, -6, 22, -21, 76, 5, 8, 5, -108, -48, 96, -92, -128, 121, 23, 31, 60, 10, -128, 8, -44, 18, 23, 10, -47, 37, 81, -106, -58, 85, 127, -95, -98, 18, 102, -52, -111, 127, 127, -81, -103, 91, 23, -100, -7, 101, -76, -81, 127, -8, -124, 127, -18, -68, 111, -37, -39, 36, 54, 13, 91, -8, -27, -38, 38, 42, -80, 87, -11, -65, 33, 60, 127, 5, -48, -45, -28, 71, 6, -85, -73, 102, -5, -81, 127, 50, -128, -70, 121, 58, -88, 12, 79, 18, -55, -55, -73, 80, -22, -74, 127, -39, -23, 93, 16, -80, -90, 38, 0, 95, 70, -103, 0, 96, -31, -29, 11, 33, 33, -87, 127, 81, -103, 27, -11, -108, -16, 92, 88, -93, 5, 39, -81, -26, -1, -33, 66, 23, -45, 57, -57, -112, 127, 54, -45, -76, 55, 101, -73, -107, 66, 21, 6, -47, -87, 24, 22, 31, -79, -3, -8, -42, 47, 86, 44, -6, 38, -64, -97, 44, 2, 21, 47, 102, 45, -8, -128, -10, 122, -48, 16, -8, -128, 75, -45, -28, 49, 6, -28, 1, -27, -28, 95, -11, -121, 22, 11, 96, 71, -116, -57, 108, 42, -39, 31, -26, -18, 55, 97, -96, -107, 127, 71, -113, 3, 78, -128, -79, 118, 15, -128, 100, 123, -68, -111, 53, -75, -66, 119, 6, -45, 29, -63, -121, 18, 127, -31, -29, 24, -69, 71, 54, -122, 29, -3, -86, 119, 18, -29, 17, 66, -6, -78, 75, -43, 7, 78, -90, -68, 63, -50, 81, 42, -85, -68, 93, 31, -68, 31, 66, 16, -95, -11, 95, 49, -68, -1, -27, 3, -64, 22, 39, -38, -68, -38, 127, -92, -96, 76, 16, 80, -3, -76, -11, 109, -8, -117, 5, 119, 29, 42, -59, -10, -1, 64, 7, -37, 50, -128, 15, -2, 65, 3, -10, -32, -2, 93, -114, 55, -48, -44, 108, -43, 12, 64, -112, -112, -21, 70, 123, -21, -86, 114, -64, -54, 127, -24, -106, 42, 37, -128, 71, 73, -103, 28, 70, -118, -12, 7, -49, 116, 76, 24, -107, -22, 122, -38, -18, 48, 21, -74, -88, -11, 48, 24, 68, -21, 50, -45, -114, 122, -8, 93, -23, -60, 91, 57, -22, -128, 97, 60, -57, 0, -48, 33, 112, -124, -122, 122, 101, 13, -5, 2, -128, -69, 58, 70, 42, -108, 55, 64, -37, 34, -39, -8, -55, 79, 15, -48, -70, -21, 43, 47, 92, -34, -96, 66, 37, -80, -7, 23, -13, 16, 37, -10, 60, 44, 49, -93, -10, 75, 1, -59, -23, -6, 107, 54, -127, 6, 37, -18, 100, 29, 16, -5, 26, 76, -128, -49, 27, 29, 90, -37, 15, 96, -59, -98, 26, 21, -13, 127, 44, -22, -128, 52, 106, -53, -90, 31, -78, -39, 127, -29, -18, -32, 13, -3, -112, 74, 60, -116, -70, 13, 43, 80, -87, -128, 12, 118, 3, -31, 49, 101, -87, -48, 122, 49, -113, -103, 113, -12, -7, 39, 6, -37, -128, 73, -31, -39, 118, -107, -106, 57, 87, 73, -78, 31, 76, -97, -48, 113, 6, -29, 15, -26, -90, 1, 53, -23, 33, -50, 12, 15, -128, 73, -11, -74, 96, -12, -128, 57, 78, -117, 86, -31, 8, -24, 29, 54, -91, -27, 12, 127, -91, -107, 127, -1, 29, -24, 24, 33, -45, 28, -86, -128, 113, 78, -78, 8, -68, 12, 15, 21, 52, -118, 39, 29, -113, 59, -69, 15, -17, -24, 119, -100, 23, 39, -48, 23, 47, -33, -75, 52, 3, 13, 49, -79, -21, 2, 108, 24, -13, -53, -69, 69, 26, -58, -33, -33, 11, 73, 97, -58, 37, 17, -107, 31, 68, 0, -128, 1, -1, -21, 2, 33, -37, 64, 90, -91, -111, 80, -32, 73, -24, -70, 112, 10, 3, 23, -32, -128, -15, 95, -22, -8, -43, 90, -7, -111, 122, 24, 5, 66, -5, -128, -11, -11, 96, 23, -70, -23, -49, 114, -3, -44, 10, 118, 102, -15, -33, -66, 42, -81, -108, 50, 86, -15, -78, 107, 8, 11, -44, -98, 127, -38, -65, 66, -21, -1, 101, 42, -78, 39, -39, -50, 127, -60, -112, 119, -44, 50, 18, -128, 0, 90, 27, 32, 42, -59, -36, -63, -15, 96, -23, -81, -79, 107, 100, -128, -71, 65, 108, -15, -91, -48, -15, 50, 66, 6, -48, 74, 27, -17, 71, -1, -107, -13, 63, 114, 59, -128, -63, 96, -65, 88, 127, -128, 16, 93, -112, 79, -37, -119, 96, 45, -52, 27, 66, -15, 3, 5, -119, -80, 38, -34, 95, 48, -80, -18, 47, 8, -13, 98, 53, -91, 8, 47, -48, -2, -15, 57, 24, -44, 74, 69, -7, -128, -17, 90, 26, -44, -38, -59, 49, 116, -128, -32, 27, -11, 60, 22, -33, 34, -54, -96, -22, 127, 65, -103, -70, 102, -75, -12, 24, 28, 44, -128, 93, -26, -16, 88, -38, -88, 57, 0, -109, -38, 127, 33, -81, 28, -55, -64, 75, 64, -45, 21, 16, -93, -49, 127, -44, -96, 100, 11, -75, -11, 92, -34, -6, 43, 85, -76, -12, 111, -66, 11, 38, -98, -66, 7, -57, 53, 57, -12, -58, -102, 59, -29, -16, 127, -106, -10, 16, 24, -28, -27, -16, 71, 71, -54, -60, 17, 64, 59, -68, -117, 127, -16, -16, 5, 22, -86, -75, 113, 76, -18, -18, -59, 0, -49, -50, -52, -49, 127, 88, -112, -80, 122, -69, 21, 33, -100, 29, -36, -7, 127, -17, -79, 6, -3, 123, -22, -58, 15, 121, -11, 26, 68, -39, 15, -117, -59, 127, -31, -116, 93, 54, -59, -3, 36, -49, -107, -31, 127, -27, -70, 100, -13, -15, 54, -28, -91, 64, 47, -106, -12, 87, -88, -80, 97, -60, 0, 5, -75, 127, 3, -13, 22, -2, -29, -74, -22, 39, 27, -81, 64, -52, -118, 80, 109, 50, 18, -128, 1, 98, -65, -43, 27, 43, 11, -93, 33, -17, -55, -52, -8, 127, 45, -16, -32, -98, -39, -24, -26, 0, 91, -12, -43, 108, 13, 54, -16, -101, 117, -47, -128, 80, 87, 24, -71, -15, -13, -27, 127, 43, -112, -45, 74, -11, -31, 52, 65, 42, -23, 7, 29, -128, 24, 123, -54, -128, 63, -39, -37, 127, -76, -18, -8, 59, -26, -49, 11, -31, 78, -44, -102, -1, 87, 88, -65, 23, 108, -10, -111, -29, 48, -69, 34, 43, -81, 11, 106, -70, 1, 34, 66, 58, -15, -121, 3, -10, 26, -34, -10, 73, -69, 22, 18, 6, -88, 5, 18, -116, 26, 87, -10, -122, -97, 54, 98, -64, 34, 5, -81, 5, 71, -26, -69, 88, 28, 48, 45, -119, -101, 88, -33, 26, 57, 16, 2, 0, 11, -113, -60, 70, 5, -63, 127, 22, -37, 24, 8, -33, 42, 60, -58, -60, -100, 90, -24, -37, 107, 29, -22, -24, -79, -5, -6, -128, 63, 3, 42, 23, -75, -50, 106, 65, -128, 32, 121, -27, -128, 13, -8, -65, 88, 108, -11, -43, 0, 12, -93, -28, 97, -85, -22, 48, -58, -21, 69, 119, -47, -66, 7, 74, 15, -86, 5, 68, 81, -71, -74, -23, 121, 28, -121, 29, 1, 86, -43, -128, 127, 38, -27, 7, 6, -85, 68, 85, -128, -37, 66, 13, 8, 43, -87, -88, -8, 97, 96, 18, 13, -128, -119, 127, 50, -106, -21, 106, -49, -33, -38, -54, 36, 108, 68, -6, 12, -38, -58, 75, 54, -128, -22, 97, 29, 5, -43, 8, -74, -63, 81, -48, -42, 100, -80, -107, 26, 95, -52, 5, 28, -81, 87, 12, 13, -22, -109, 59, 116, -32, -60, 34, -2, -116, -3, 57, 90, -78, -66, 45, 54, -34, 27, 2, -71, -22, 74, 68, 17, 10, -101, -65, -17, -3, 124, 111, -78, 3, -6, -78, 23, -36, -11, 29, 24, 98, 55, -85, 49, 127, -69, -70, -24, -8, 109, 16, -64, 5, -26, 6, 26, 48, 54, -44, 33, -16, 97, 92, -44, -87, -102, 8, 53, 0, -11, 48, 65, 12, -44, -60, 24, -81, 43, 116, -124, -24, -1, 8, 95, -80, 6, -74, 17, 31, -88, 22, 44, 0, -22, 29, 90, -8, 8, -53, 18, 127, -36, -92, 32, -49, 44, 5, -101, 76, -33, -5, 0, -5, -6, -38, -34, 10, 60, 98, -8, -34, -76, 65, 98, -128, -80, 52, 57, 43, -31, -100, 60, -36, 6, 42, -54, 42, -109, 60, 68, -113, 23, 100, -128, -118, 92, 12, 6, 102, 80, -11, -112, -111, 106, -1, -42, -26, 80, -15, 47, 16, -85, 76, 11, -87, -15, -11, 127, 11, -128, 65, 97, 11, -52, 0, 29, -11, 2, -128, -23, 117, 24, 0, -128, 15, 27, -55, 103, 57, -81, -26, -58, 50, 0, -15, -65, -5, 127, -128, -109, 11, 113, 102, -5, -117, -10, 75, -97, 2, 114, 12, -76, 24, 43, -70, -10, 81, 28, -107, 24, -1, -101, -1, 59, 75, 97, -36, -108, 90, 29, -102, 70, -32, -114, 96, 26, 10, -45, -16, -15, 100, -34, -63, 93, 17, 21, -116, -12, 80, -22, -37, 90, 10, -71, -48, 127, -6, -53, 21, -52, 6, 97, 127, -76, -26, 29, 0, -47, 15, -48, -32, 85, -52, -107, 42, -2, 92, 39, -47, -23, 48, 69, -128, -53, 26, 15, 32, 29, 97, 2, -53, 73, 90, -98, -119, 93, 111, 15, -128, 10, 0, 12, 43, -43, 42, 32, -57, -42, -38, -73, 127, -42, 5, 127, -128, 22, -48, -63, 21, 57, 75, -64, -45, 28, 34, -29, -75, 29, 16, -28, -10, 47, -47, 64, -26, 26, 65, -52, -26, -128, 92, 50, -128, 88, 27, -69, 57, -10, 22, -119, -68, 127, -3, 21, -37, -86, 22, 64, 58, 7, -128, -64, 88, 7, -52, 93, 2, 44, 7, -12, 71, -98, -75, -15, 0, 127, 48, -128, 1, 103, -81, 69, 15, -34, 57, -11, 34, -117, -63, 127, 69, -91, 31, -39, -29, -52, 60, 108, -37, -107, -18, 64, -5, -128, 57, 127, -52, -91, 38, -59, -122, 8, 16, 70, 90, 45, -118, -10, 127, -44, -80, 59, 81, -101, 52, 21, -123, 103, -5, -111, 7, 127, 69, -49, -6, -49, -34, -6, -111, 34, -57, -54, 127, -92, 5, 50, -13, 43, -128, -1, 29, -39, 6, 123, 13, -128, 8, 90, 79, -47, -31, -90, -10, 91, -108, 12, 49, 53, -47, -27, 58, -73, -93, 63, 53, -119, -21, 70, 101, -43, -128, -2, 114, 12, -76, -6, 71, 45, 50, -23, -116, 50, 63, 8, -76, 6, -7, 2, 29, -23, -33, -45, -65, 69, -13, -128, -16, 127, 57, -114, -38, 127, -2, 42, -55, -28, 3, 47, -12, 87, -8, -97, 108, 85, -98, -107, 123, 69, 31, -44, -68, 48, -80, 63, 66, -87, 50, 16, -123, -26, 100, -26, -96, -16, 47, 23, 66, 0, 38, 43, -112, 60, 80, -34, -52, 12, 12, -128, -29, 75, 3, 34, -92, -23, 68, 5, -121, -15, 53, -45, -71, -1, 124, -53, -50, -24, 21, -13, 3, 28, 37, 49, -108, 5, 44, 37, -11, -76, -57, 127, 116, -85, -6, -92, -54, 93, -75, 21, 23, 8, -53, -16, -2, -65, -18, -43, 86, 117, -90, -87, 8, 127, 76, -128, -22, 6, -59, 127, 44, -128, 100, 24, -13, 38, -34, -80, -2, -58, -27, 52, -38, 116, -15, -8, 17, -24, 80, 71, -109, 23, 122, -128, -3, 63, -39, -79, 80, 54, -128, -7, 102, 78, -12, -90, 3, -16, 26, -49, -45, -31, 12, 70, -128, 48, 28, -87, -7, 122, 123, -128, -32, 109, -57, -68, 15, 98, -12, -100, 17, 48, 27, -75, 11, 44, 31, -34, 57, 27, -53, -17, 27, -50, -106, 111, -54, -43, -6, -31, 66, -38, 38, -17, 78, 117, -118, -81, 79, 66, -47, -98, 0, 10, 1, 127, 3, 22, -85, -52, 81, 58, -103, -24, 37, -8, 32, 12, -86, 36, 117, -70, -13, -39, -34, 53, -80, 43, 86, -31, -65, -75, -76, -54, 113, 37, 42, -59, -71, 127, 1, -21, 15, -48, -55, -79, -5, -12, 111, 23, -8, 49, -128, 27, 18, 0, 28, -29, 33, -17, -8, -21, 80, 27, -109, -3, 118, -97, -32, 34, -75, 18, 23, 127, -79, -1, 26, -74, 127, -80, 0, 100, -18, -3, -69, -116, 26, 127, -8, -128, 1, 11, 38, 29, 49, 66, -3, -28, 22, -68, 15, 79, -78, -128, 85, 37, -2, -109, 13, 107, -128, 5, 69, -128, 32, 8, -65, 127, 95, -87, -128, -36, 124, 15, -36, -1, -31, -8, 127, 106, -111, -13, 70, -128, 45, 102, -88, 11, 23, -81, -16, -81, -45, 60, -33, 101, 18, -112, 100, -18, 0, 75, -90, -52, -43, 70, 58, -107, -117, 91, 29, -28, 44, -53, 31, 37, 79, -66, -85, 127, 48, -128, 85, -27, -59, 16, 81, 96, -124, 5, -38, -71, 93, 48, 10, -128, 3, 102, -76, 22, -26, 5, -36, 28, 88, -34, -109, 31, 96, -57, -29, 7, 5, 0, 10, -86, 49, 63, 39, -86, -65, 31, 39, -24, 113, 18, -128, 86, 127, -63, -90, -7, -24, 50, 127, 29, -128, -90, 93, 112, -10, -128, 3, 24, 42, 127, -92, -86, 58, 127, -54, -37, -17, 16, 93, -124, 68, 87, -70, 22, -92, -108, 24, 58, 78, -36, -45, 116, -10, 15, 27, 7, 15, -17, 22, -119, -23, 127, -88, 3, 79, -92, -43, -73, -22, 58, 0, -6, 127, 86, -128, -70, 127, -42, -42, 54, -47, 68, -47, -6, 52, 10, -8, -65, 44, 23, -6, 127, -64, -43, 127, 47, -128, -71, 127, -54, -44, -26, -10, 79, 69, -55, -21, 47, -45, -74, -52, 103, 108, -128, -79, 24, 76, 23, -70, -75, 79, 55, 27, 3, -128, 42, 85, -113, -60, 100, 29, 7, 21, 8, -88, -23, 5, -78, 33, 127, -38, -49, 63, -66, 36, -69, -8, 81, -12, -113, 36, 32, -23, 54, -118, 29, 44, -2, -113, 12, 65, -50, 11, -47, -8, 101, 43, -34, -128, -36, 127, -15, 47, -23, -31, 52, -63, -52, 0, -45, 32, -13, 17, -1, -96, -45, 38, 127, 65, -103, -36, -3, 63, -75, -21, 43, -111, 74, 17, -88, 127, 98, -116, 22, -38, -96, 108, -91, 49, 54, -107, 52, 71, -97, -85, 6, 32, 69, 102, -98, 16, 33, -70, 49, -10, -102, -63, 98, -79, -33, 127, 39, -113, -86, 95, 26, -44, -16, -12, -3, -97, -66, 78, -13, 12, 109, -58, 36, 1, -92, 127, -32, -26, 74, -119, 15, -15, 15, 59, -65, -27, 70, 5, 36, 101, 68, -114, -58, 85, 70, -117, 16, -27, -27, 127, -44, -96, -34, 22, 85, 6, -37, 80, 117, -13, -47, -65, 18, -60, 5, 90, -121, -100, -38, 116, 114, -22, -7, -122, -52, 95, -38, -88, 98, -76, -86, 85, 3, -5, 54, 54, -28, 6, -38, -26, 43, -53, -59, 73, 80, -86, 6, 127, -70, -63, 98, -70, -32, 101, -13, 47, -23, -1, -49, -60, -49, 42, 127, -97, 26, 15, -128, 48, 32, -16, 127, 23, -81, -101, -15, 28, -7, 108, 127, -91, -128, 101, 36, -32, -16, 74, -15, -10, 39, -33, -106, 22, -2, -103, -23, 33, 91, -65, 31, 92, -95, -7, 1, -127, -98, 127, 18, -128, 93, 21, -29, 74, 70, -3, -128, -60, 101, 47, -106, 6, 43, -11, -1, -93, -81, 127, 54, -23, -91, -27, 98, 11, -66, -33, -80, 31, 76, -50, 49, -47, 1, 127, -2, -106, 34, -108, 29, 87, -28, -86, -42, 45, 101, -96, -36, 127, 23, -128, 13, -34, 10, 60, 7, -65, -128, 127, 80, -80, -103, -2, 69, 32, -45, -48, -17, 0, 39, -39, 118, -17, -96, 44, 57, -24, -18, 10, -6, 34, 49, -44, 29, 28, 48, 6, -23, 76, -65, -57, 26, 7, 74, -102, -73, 59, 26, 21, 28, -128, 31, 117, -118, -73, 5, 127, 13, -44, -48, 38, 124, -50, -13, -42, 31, 1, -2, -2, -55, -37, 117, 86, -60, -6, 34, -128, -81, 93, 73, -106, -5, 74, 21, 10, -50, 16, -26, -128, 2, 100, 23, -69, -64, 38, 64, 79, 10, -116, -58, 127, -17, -128, 123, -49, 48, 108, -128, -43, 44, 108, -33, 6, 3, -128, 70, -15, -78, 53, 10, 59, -64, 65, 127, -128, -70, 74, -48, 117, 73, -128, 70, 87, -127, -22, 88, -87, -50, -44, 47, 127, -128, -102, 127, 45, -95, 17, 60, -15, -124, -39, 74, 7, -6, 44, 44, 34, 68, -12, -24, 5, 65, -3, 103, 75, -59, 13, -124, -58, -17, 121, 13, -123, 6, 24, 122, 27, 11, -12, 43, 22, -87, -79, 63, 39, -88, 76, 45, -29, -128, 52, 112, -101, -128, 101, 6, 6, 63, -87, -85, 74, 0, -57, 88, -42, -42, 10, 36, -59, 28, 48, -5, -90, 0, 24, -15, -98, -32, 81, -118, 29, 81, 24, -101, -15, 95, -64, -17, 1, 45, 32, -121, -66, 27, -22, 66, 100, -39, -71, -74, 38, 7, -49, -16, 17, 127, 80, -111, -55, 27, -8, -57, -23, 47, 16, 96, -75, 5, 45, -43, 39, -55, -112, -13, 127, -17, 21, 49, -8, -80, 5, 0, -42, -74, -6, 127, -121, -39, 52, 18, -65, 53, 98, -122, -74, 0, 5, 45, -45, 80, -6, -128, 55, 58, -17, -13, 92, -28, 66, 52, -78, 60, -81, -69, -1, 108, 8, -92, 33, 95, -103, 0, 119, 26, -128, -92, 57, 49, 69, -18, -44, -71, 37, 127, -65, 7, -66, -109, 127, 116, -88, -78, 42, 26, -12, -128, 17, 27, -52, 18, -32, 42, 127, 53, -109, -112, -5, 127, 52, 31, -70, -128, 127, 80, -33, -86, -45, 97, -57, -66, 98, -95, -116, 127, 109, -12, -37, -49, -100, -58, 127, -16, -48, 107, -98, 39, 109, -128, -8, 24, 95, 33, -128, 74, 0, -117, 0, 127, -70, -24, 53, 37, 13, -92, 11, 8, -52, 3, -28, 23, 58, 65, -2, -128, 34, 96, 11, -74, 10, -28, -17, 74, 13, 2, -47, -98, -80, 127, 1, -122, 95, 65, 71, -90, -128, 116, 98, -55, -98, 98, 103, -69, -11, -34, -13, -7, -75, 27, 95, 49, -32, -101, 8, 33, -66, -26, 113, -11, -95, 127, 1, -31, 33, -59, 76, 8, 23, -22, -15, 81, -122, -27, 44, 64, -95, -107, 87, 5, 55, -15, -57, 54, 57, 65, 37, -37, 28, -47, -18, 91, -121, 32, 27, -52, -36, -50, 127, 101, -106, -37, 47, -7, -97, -42, 88, -12, -33, 122, -38, 11, -93, -45, 36, -2, -8, 86, 93, -11, -128, -42, 109, -58, -38, -17, 85, 37, -102, 60, 2, 10, -6, -86, 33, 73, 7, -97, 90, 127, -128, -64, 127, -90, 24, -8, -59, 127, 44, -128, 22, -60, 10, 80, -90, -58, 93, -34, 8, -39, 55, -17, 2, 16, -71, 5, 101, 71, -123, 12, 66, -76, -81, 85, 29, 55, 22, -39, 28, -45, -128, 64, 68, 11, -52, -128, 5, 49, 3, 127, -21, -116, -3, 11, 79, 37, -12, 2, -24, 59, 127, -8, -47, 36, -103, -128, 127, 96, -36, -42, -64, -119, 50, 13, 70, 113, -128, -100, 26, 71, -22, 15, 92, -78, 16, -26, 11, -27, -12, 123, 1, -59, -1, 5, -11, 70, 8, -86, 52, 3, 69, -64, -81, 91, -16, -21, 47, 28, -6, 42, -97, 21, 27, 26, -66, -112, 127, 58, -128, 6, 47, 29, 59, -6, 24, -128, -49, 66, -15, -49, 103, 22, -81, -10, 123, 33, -64, -6, -50, -18, 45, 28, 117, 42, -128, 79, 88, -128, 3, 116, -21, 18, -31, -74, 65, 3, -26, 127, 17, -52, -96, -11, 127, -64, -54, 92, 22, -128, -71, 127, -34, -76, 127, 49, -65, 13, -45, -114, 91, -95, 32, 36, -42, -29, -5, -7, -13, 123, -75, -111, 102, 5, 11, 49, -27, 114, -54, -128, 127, -12, -22, 114, -101, -31, 49, -116, 12, 12, -29, 52, -49, -7, -44, -59, 127, 63, -100, -53, 50, 22, -28, -65, 58, 119, -68, 21, 34, -92, 37, -1, -52, 5, -22, -102, 5, 36, -18, -31, 80, -59, -114, 63, 108, -44, -28, 68, -117, 68, 127, -97, -86, -34, 55, -55, -50, 42, -23, 127, 63, -15, -17, -106, 42, -31, -7, -3, 36, -58, -3, 87, -90, -128, 12, 48, 2, 119, -101, -60, 127, 58, -128, -63, 54, 65, -3, -48, 75, -38, -64, 24, -3, -52, -47, 47, 93, 57, 10, -47, -116, 57, 48, -26, 43, 8, 11, -128, -5, 111, -57, -45, 32, -6, -128, -47, 90, 29, 37, -31, -124, 24, 2, 48, 88, -96, 86, -15, 13, 64, -53, 55, -74, -119, 80, -18, 88, 39, -121, 71, -5, 39, -3, -109, 65, 29, -21, -43, -52, 48, 102, -60, 22, 73, -23, -87, 29, 28, -71, 33, -38, -73, 101, 60, -57, -36, 93, 0, 13, 109, 18, -1, -27, -98, -57, 47, 109, 34, -47, 45, -92, -80, 127, 45, -37, -18, -128, 43, 21, -28, 24, -8, 32, 73, 22, -55, 26, -80, -3, 8, 57, -13, 38, 0, -81, -49, 78, -3, 15, 0, 50, 59, -113, 55, -7, -100, 45, 12, 58, 13, -24, -93, -108, 37, 127, 28, -48, -12, 0, -86, 27, 24, -69, 55, -111, -122, 127, 85, -128, 1, 127, -116, -71, 53, 118, 32, -76, -11, -66, 33, 11, 85, 55, -127, -54, 78, 101, 29, -128, -13, -1, -73, 21, 127, -69, -76, 127, -85, -109, 34, 96, 127, -128, 10, -2, 37, 12, -48, -5, -22, -44, 36, 29, 18, 47, -54, -76, 32, 5, -11, -32, 34, -118, 18, 127, -128, -68, 127, -42, -60, 121, 39, -119, 39, 21, -91, 66, -100, -87, 70, 53, 2, -90, -29, 54, 127, 27, -53, -6, -79, -12, -7, -33, 65, -18, -58, 108, 47, -128, 96, 119, -50, -38, -114, 38, -6, -5, 54, -74, -103, -7, 8, 76, 16, -50, -43, 38, 7, 100, -18, -38, 54, -17, 81, -100, 12, -6, 38, 27, -118, 127, -7, 48, 32, -90, 57, 57, -107, -21, 12, -11, -80, 54, 33, -31, -26, 0, 127, -48, -98, 127, 45, -74, -39, -5, 45, -79, 15, 53, -39, 54, -38, 3, 73, 3, 69, -65, -50, -5, 90, 75, -48, -128, 16, 13, -23, 107, -15, -79, 88, 42, -123, 17, 0, 32, -37, 54, 88, -52, -88, 100, -28, -97, 71, 54, 64, -75, 39, -18, -49, 121, -78, -68, 127, 52, -85, -73, 23, 98, -16, -87, 3, 55, 47, -26, -108, 59, -2, 11, -23, -59, 80, -42, 0, -64, 64, 31, -109, 74, 22, -2, -23, -3, -80, -31, 79, 10, 8, 71, -66, -122, 15, 116, 69, -128, -26, -5, 103, 87, -24, -98, -90, 87, 36, 24, -7, -74, -57, -64, 8, 127, 45, -45, -59, 15, -88, -116, 58, 119, -96, 23, -33, -47, 108, 45, -24, -128, 92, 45, -18, 33, -21, -119, -12, 68, -63, 8, 2, 55, 58, -16, 21, -8, -10, -6, 16, 76, -7, 44, -1, -50, 36, -24, 55, -52, -93, 60, 7, -53, 127, -43, 11, 87, -128, -10, 0, 2, 113, -48, 49, -26, -13, 38, -26, 109, -18, -18, -11, 23, -5, 16, -36, -103, 44, 28, 18, 65, 38, -2, 0, -17, 5, 1, -90, 71, 106, -121, -102, 80, 27, 60, 1, 2, -96, 27, 78, -85, -23, 98, -91, 1, 86, -118, 53, -90, -34, 44, 6, -27, 73, -23, -16, 48, -11, 49, -76, -42, 127, -64, 7, -18, -117, 60, -7, -12, 36, 80, 37, -16, -16, 0, -26, -68, -66, 37, 17, 31, -116, -90, 34, 127, 0, -11, -12, 39, 5, -58, -10, -22, 96, -54, -11, -52, 15, 116, -97, -123, 81, -5, -109, 96, 2, 63, -23, -31, 70, 24, -29, -32, 71, -26, -74, -39, -7, 111, -50, 28, 18, -31, -3, -39, 127, -68, -60, 127, -111, 59, -34, 3, 22, -114, 69, 34, 85, -6, -5, -21, -96, 13, -22, -12, 127, 15, -87, -18, -7, 58, 123, -18, -128, -15, 127, -69, -52, 65, 78, -5, -93, 95, -32, -58, 117, -13, -33, 22, -128, 11, 11, -34, -23, 0, 87, 90, -15, -8, -128, 27, 37, -128, 38, 66, -18, -21, 27, 60, 12, -70, -57, -27, 33, 87, 48, -47, -43, 65, -12, 16, 26, 7, 118, -49, -2, 27, -74, 32, 27, -5, 7, 75, -8, 16, -54, 21, -33, 2, 52, 8, -98, 3, 118, -96, -87, 29, 53, -13, 45, 7, -28, 39, 6, -88, -124, 33, 117, -63, -128, 7, 127, -5, 53, -58, -102, 29, 127, -1, -128, 76, 38, -65, 50, 1, 34, 79, 1, -88, -49, 76, 100, 55, -78, -8, 0, -3, -5, -39, 127, -18, -63, 58, 24, -39, 10, 58, -42, -26, -76, 11, -1, -26, 81, -1, -34, -57, -36, -2, 31, 26, 43, -45, -52, 127, 58, -85, -38, 85, 29, -111, -50, 0, 127, 90, -73, -37, 32, -63, -53, 127, 64, -87, -70, 31, -36, -75, -15, 102, 33, -34, 98, 47, -114, 33, 31, -128, -17, 127, 28, -17, -128, 28, -29, -128, 127, 74, -48, -33, 43, 53, -100, -6, -1, 26, -26, -7, -79, -10, 63, -34, 109, -36, -102, 47, 6, 108, -7, -42, 100, -93, -28, 127, -116, -48, 127, 5, -128, -13, 22, -75, 49, 101, 29, 15, -48, -109, 37, 47, -5, 49, 1, -74, -123, 97, 88, -128, 27, -53, 29, 74, -117, -8, 76, -32, 76, 27, -128, -21, 24, 55, 15, 42, -38, 101, 26, -57, -39, 97, -42, -15, 117, -7, -122, 23, 78, -128, -70, 117, -23, -70, 34, 55, 32, 60, 12, -65, -44, 68, 26, -50, -70, 73, 127, -128, -2, 16, -1, 91, -103, 6, 64, -124, 29, 127, -128, -26, 5, -3, 36, -7, 59, 18, 16, 85, -95, -85, 47, 36, 101, 22, -24, -128, -16, 127, -93, -50, -6, 123, -11, -78, 98, 63, -45, -69, 69, 18, 17, 23, -13, 24, 5, -128, -68, 74, -36, 12, 107, -39, 39, 28, -128, 45, 57, -13, -38, 16, -98, -13, 109, -101, 60, -8, 12, -15, -47, 52, 34, -58, 108, -8, -2, 80, -111, -81, 0, 49, 66, -112, 59, 75, -50, -81, -10, 37, 78, 85, -128, 31, 36, -22, -78, -55, 127, 48, -103, -57, -33, 127, 16, -124, 3, 44, 127, 7, -68, -39, -55, 29, 43, -47, 119, 127, -128, -69, 31, 127, -37, -100, 127, 29, -128, 65, 109, -17, -60, -111, -45, 101, -32, -17, 114, -79, 15, 50, -17, -63, -128, -44, 127, 31, -123, 87, 24, -88, 127, 24, -128, -42, 127, -44, -1, 127, -10, -69, -7, -39, 17, -87, -74, 16, 93, -12, -29, 76, 68, -59, -121, -26, 71, 127, -45, -60, 27, 8, 6, -37, -78, -91, 117, 11, -106, 106, -18, 102, -15, 2, 50, -128, -50, 127, 0, -10, 108, -42, -111, 60, -71, -32, -16, 29, 74, -32, -39, -32, 28, -22, 107, 64, -128, 23, 108, -93, -91, 127, -21, -76, 113, 38, -74, 28, -3, -22, 7, -32, -12, -70, 37, 92, 8, -8, -53, -28, -10, 81, 52, -33, 48, -17, -106, 123, -47, 32, 0, -107, 127, -11, -26, 34, 58, 54, -128, -59, 60, 52, 21, -2, -27, -118, -27, 12, 50, 32, -68, 28, -60, -128, 47, -2, 28, 55, 68, -27, -87, -68, 85, 2, -48, 26, 70, -1, -74, 127, 52, -44, 11, -39, 3, -5, 38, -74, 37, 58, -10, -38, -45, -42, 27, -50, -12, 24, 34, 23, 28, -81, -12, 80, -69, 71, 54, -28, 38, -29, -69, -21, -22, -45, 114, 96, -81, -43, 73, -53, -119, 114, -81, 29, 18, -22, -50, 16, 127, -47, -128, 31, 66, -12, -106, 49, 26, -17, 8, -68, -16, 118, 23, -70, -106, 23, 55, 10, -50, -5, -11, 26, 55, -63, 26, 87, 49, -55, -73, 73, -73, -10, 53, 23, -55, -18, 43, 0, -48, -79, -34, 127, -13, 18, 28, -88, 12, 96, 57, -68, -87, -68, -10, 127, -15, -15, 55, -80, -42, 127, 108, -128, -27, 45, -92, 113, -26, -15, 85, -65, 37, 16, -111, -92, 68, 96, -64, 50, 13, -121, 11, 106, -73, -28, 53, -36, -55, -44, 79, 34, -81, 50, 87, 3, 44, -15, -58, -96, 17, 33, 34, 3, 60, 59, -117, -45, 21, 37, -26, -101, -28, 16, 13, 74, 102, 15, 5, 13, -38, -92, -86, 75, 73, -29, -97, 3, 3, -128, 86, 127, -128, -54, 28, -28, 15, 90, 38, 5, -48, -101, -63, 97, 29, -78, -5, -2, 127, -29, -124, 127, 54, -73, 24, 13, -52, -39, 28, 127, -50, -81, 127, 2, -2, -54, 6, 127, 2, -128, 37, -13, -33, -54, -52, 27, 42, 57, -5, 0, 57, 5, 96, 80, -78, -55, -38, 66, 15, -39, 0, -2, 31, -64, -116, 59, 55, 26, 8, -74, 116, -2, -58, 48, -47, 23, 24, -36, 49, -11, -47, -91, 45, 37, -128, 18, -7, 13, 34, 38, -57, 65, 3, 5, -29, -78, 33, 36, 81, -6, -47, 21, -127, -53, 79, 24, -60, -28, 38, 0, 127, 108, -122, 3, 8, -45, -27, 31, -63, 37, 39, -90, 73, 76, -116, 53, 127, -112, -86, 102, -66, -102, 127, -13, -21, -3, 39, 52, -87, 49, 39, -128, 42, -27, -93, 63, 102, -5, 43, 27, -128, -49, 127, 44, -24, 10, -76, -5, -47, -128, 107, 60, -98, 21, 76, 15, -12, -57, -44, -48, 23, 6, 21, 13, -8, 64, 24, 59, 48, -109, -24, -63, 37, 58, 11, 2, -65, -12, 6, 63, -8, -81, -10, 91, 52, 36, -70, -75, 10, 59, -8, 2, -109, -102, 48, 57, 75, 43, -57, -8, 127, 29, -106, -6, -23, -38, 5, 88, 60, -16, -47, 85, 33, -90, -2, -26, 0, -63, 95, -39, 29, 53, -27, 55, -101, 10, -81, 27, 22, -109, 5, 17, -45, 78, 127, -122, 7, 101, -44, -108, -29, -39, 7, 12, 68, -45, 16, 36, -76, 80, 26, -55, 0, 49, 10, 96, 8, -38, 93, 42, -12, 47, 29, -69, -50, 21, 26, -74, -11, 11, 16, -96, 2, -5, -49, 38, -18, -64, 88, 36, -34, 81, -50, -45, -64, 10, 17, -43, 107, 58, -10, -85, -7, 49, 43, -91, -63, 101, 32, -108, -22, 79, -3, -49, -59, -23, 127, 32, -121, 55, 102, 0, -57, -64, -13, 54, 60, -48, 1, -7, -106, 18, 85, 22, -128, 11, -36, 7, 60, 6, 34, 7, -90, -85, -10, 27, 26, -63, 92, 42, -37, 15, -71, -44, -36, 92, 127, -5, -128, 10, 15, -38, 1, -33, 12, 50, 95, -53, -117, 39, 3, -49, 58, 92, -17, 16, -78, 37, 111, -128, -32, 103, 8, 8, 6, -36, -75, 16, -11, -11, -1, -128, -21, 127, -49, -38, 50, -70, -60, 112, 85, -111, 49, -32, -128, 81, -3, -10, 68, 116, -59, 3, 42, -128, 66, 59, -5, -39, -57, 32, -43, 117, 16, -97, 96, 17, -128, -7, 127, -73, -96, 96, 34, -97, 73, 38, -65, 36, 16, -128, 37, 8, -128, 91, 18, 64, -47, -101, 53, 73, 47, -18, -6, 96, 38, -111, -18, 92, 16, -71, -96, -24, 32, 117, 12, -92, 42, 0, -23, 70, 23, -37, 91, 21, 1, 101, -113, -12, 127, -90, -118, 48, 88, 8, -52, -6, 98, 60, -114, 0, 21, -32, 91, 1, 52, 73, -101, -81, -60, 71, 102, -90, 24, -3, -15, 15, -58, 68, 118, 23, -52, -8, -103, -79, 29, 18, 47, -68, -52, 127, 47, -85, 87, -58, -29, 127, -121, -78, 57, -3, 108, 109, -106, -43, -31, 75, 88, -123, -32, 91, -44, -53, 92, 27, -18, 69, 37, -128, -114, 15, 127, 47, -100, 48, 38, -128, 18, 117, -106, 26, 79, -5, -42, -128, -17, 123, -96, -65, 32, 48, 127, -64, -15, 31, 13, -45, -33, 85, -16, -33, 68, -34, -101, 21, 22, 116, -2, 11, 34, -55, 27, -18, -10, -3, 15, 107, -100, -26, 7, -54, 127, 96, -128, -34, 12, -86, 96, 95, -32, -100, -53, 66, 42, -39, 34, 32, 43, 22, -128, -34, -2, 73, 58, -44, -108, -38, 93, -28, 48, 48, -97, 28, 8, -8, -57, 32, 59, -128, 11, 58, -81, 93, -93, 10, 21, -24, 32, -69, 27, 79, 7, -5, -23, -47, -17, 44, 48, -124, -98, 127, 101, -58, -38, -2, -36, 100, -1, -128, 127, -39, -42, 65, -103, 85, 24, -49, 26, 69, 13, 23, -27, -91, 48, 127, -23, 0, -5, -91, -95, 93, -12, 37, 2, -21, 2, -2, 47, 12, 18, -11, 23, -52, 64, 55, -21, 57, -24, -5, -48, -124, 48, 100, -79, -100, 91, 116, -128, -50, 55, -27, -8, 53, 127, -58, 0, 118, -73, -128, -3, 127, -26, -11, -87, -76, 74, 91, -48, -87, 116, 78, -74, -33, 43, 42, 1, -64, 22, 68, 0, 26, 7, -42, 70, -43, -48, 60, -60, -92, 111, 69, -128, -31, 90, -53, 5, 112, 3, -53, -128, 3, 55, -48, 86, 48, -15, -111, 36, -26, -8, 5, 31, -32, -3, 71, -44, -64, -1, -74, 39, 55, 5, 31, -5, -85, -128, 52, 59, -100, 7, 87, 18, 12, 26, -70, -50, 39, 15, -66, 45, -23, -29, 45, -24, -45, -15, -17, -78, -7, 85, 76, 16, -88, -3, 42, 5, -3, -103, -69, 93, 39, -128, -1, 87, 42, -103, -101, 114, 91, -31, -37, -48, -8, 18, 102, 58, -28, -93, -128, -5, 127, 78, -128, -34, 106, 53, -59, -33, -17, 68, 26, -128, 106, -26, -15, 117, -121, 37, 11, 22, -24, 3, -57, -2, 12, -92, 107, -3, -7, 87, -39, -16, 28, -28, 81, -64, -91, 53, 78, 26, -76, -28, 91, 127, -88, -103, 123, -8, 70, -63, -102, 76, 118, -24, -124, -2, 80, 97, -58, 63, -13, -47, 12, 23, 78, -122, 11, -42, -37, 59, -5, 18, 0, -92, 26, 109, -58, -68, 127, -18, -101, 17, 88, -12, 3, 98, -68, 75, -1, -75, 108, -5, 32, -76, -96, 127, -1, -114, -34, -7, 124, 73, -17, -74, 32, -22, 44, 109, -122, 0, 119, -87, -11, 8, -48, -38, 119, 17, 3, -80, -5, 79, -54, -3, 33, -128, 2, 64, -98, 81, 3, 13, -21, -128, -27, 127, -36, -13, 100, -108, -26, 63, 23, -92, 85, 112, -128, 26, 13, -107, -22, 39, -13, 119, -13, 29, 92, -43, -80, -121, 69, 121, -128, -108, 127, -29, -128, 127, 90, -68, -101, -50, 27, 100, -6, -87, 74, 49, -92, -65, 127, 0, -76, 117, -79, -38, 127, -124, -31, 64, -47, 6, 28, 12, 34, 0, 12, 54, -13, -10, 17, 60, 50, 13, -34, 75, 63, 7, -71, 2, 100, -128, -113, 74, 0, -15, 127, 86, -128, -58, 12, 0, 63, -7, -15, 66, -38, -12, -75, -23, 112, -88, -128, 27, 127, -39, -95, 53, 127, -29, -128, 127, 38, -118, -13, 70, 21, -64, 18, 69, -8, 2, -107, -59, 26, 74, -24, -128, 93, 75, -37, 5, -128, 39, -16, 8, -31, -79, 53, -22, 87, 48, -92, -7, 127, 7, 31, -47, -3, 39, -112, 37, 54, -17, -52, -53, 87, 98, -68, -15, 59, -53, 0, 91, 101, -48, -74, -65, 68, 93, -119, -22, 6, -11, 85, 85, -13, -60, -75, 11, 127, -52, -128, 76, 127, -85, -6, 12, 44, 58, -33, -92, 36, 102, -32, -38, -60, -76, 92, -23, -118, 3, 127, 2, -38, 16, 119, 79, -74, -128, -18, 114, -11, -29, -6, -22, 81, 100, -38, -48, 23, 124, -5, -128, 112, -7, 18, -1, -52, 80, -15, -34, 53, -85, -1, 127, -98, -60, 95, 24, -60, -123, 2, 123, -38, -55, 69, 31, -128, -85, 13, 66, 127, -43, -79, 68, 0, -69, -68, 0, 21, 92, 76, 22, -1, -101, 36, 98, -27, -66, 7, -57, 7, -18, -69, 0, 122, -28, -124, 127, 0, -128, 74, 18, 12, 111, 57, -128, -97, 127, -48, -107, 80, 59, 73, -128, 10, 78, -10, -24, -123, 49, -52, -85, 38, 54, 29, 109, -5, -103, 97, 26, -90, -45, 76, 80, -128, 0, 117, -97, -8, -66, 15, 17, 23, 57, -90, 24, 0, -47, 7, 75, -49, -32, 127, -60, 11, -17, -66, 37, 53, 127, 11, -44, -79, -23, 68, -17, -53, 26, 85, 49, -70, -76, -45, 3, -7, 42, 127, -58, -15, -24, -119, 127, 55, -22, -107, -65, 127, -58, -58, 32, -29, 3, 0, 65, 96, 13, 16, 29, -128, -12, 113, -7, -122, -68, 26, 45, 111, -48, 37, 60, -63, 75, -2, -121, 85, 66, -52, 21, 37, 23, 2, -22, -2, -6, -128, -21, 37, 80, -43, -64, 57, -66, -42, 113, -18, -68, 127, 57, -128, -10, -13, 27, 11, -7, 42, 44, 27, -18, -111, -48, 54, -74, -39, 85, -71, 23, 8, -1, 73, -2, -76, -23, 127, -5, 36, 76, -85, -12, 0, 6, -75, 13, 2, -31, -3, -90, 65, 32, 68, 69, -45, -53, -121, -32, 38, -13, 106, -2, -27, -17, 24, 28, -73, -22, -91, 13, 64, 22, -28, -71, 59, 71, 55, 32, -128, -80, 127, 43, -78, 31, 0, -71, -10, 54, 7, -1, -128, 0, 24, 32, -49, -86, 95, 52, 6, -27, -109, -44, 24, 37, -1, 54, -65, -58, 119, -24, -3, 42, 69, -95, -59, 100, 10, 63, -43, -95, 92, 16, -128, -16, 80, 0, 32, -22, -60, 70, 127, -55, -3, -45, 33, -37, 17, 106, -128, -37, -55, 86, -27, -128, 127, 26, -74, 22, -44, 79, 63, -128, -36, 127, -33, -128, 17, 28, 1, 71, 69, -70, 68, 32, -86, 71, 24, -76, 39, -70, 60, 100, -15, -128, 7, 127, -108, -75, 7, 66, -26, -86, 113, 71, -128, -55, 117, -13, -57, -79, 109, -18, -119, 127, 22, -48, 18, -87, 93, 7, -127, 127, -26, -111, 127, 117, -128, -64, 73, 39, -48, 55, 113, -128, 13, -2, 5, 78, 11, -81, 29, 91, -93, 66, 17, -17, -12, 48, 50, -119, -76, 127, 127, -128, 5, 100, -7, -2, -128, -49, 68, -33, 127, -34, -118, 124, -28, 45, -13, 13, 98, -15, -92, 55, 17, -42, 7, 36, -23, 70, 53, -128, 17, 58, -70, -6, 22, -26, 0, 37, 36, 16, -6, -17, 10, 31, -113, 33, 45, -97, 16, 127, 22, -107, 13, 71, -11, -7, -68, -128, 116, -2, -87, 80, 66, 0, -123, -44, 127, -7, -37, 8, 59, -75, 22, 39, -32, 65, -123, -122, 127, 29, -128, 53, 123, -13, -71, -2, 7, 37, -16, -74, -100, 116, -45, -1, 81, -128, -55, 97, 50, 17, 75, -87, -3, 66, -13, -48, -22, 59, -33, -53, -44, 17, -29, -55, 34, 74, 75, -128, -1, 88, -52, 33, -15, -45, 21, -90, 12, 78, -22, -113, -15, 86, 0, -50, 15, 13, 76, 127, -122, -71, 107, 10, 60, 23, -55, -79, -15, 49, -34, -48, 2, -36, -3, 127, 29, -13, -101, -70, 96, 53, -68, 48, -58, -15, -33, -31, 127, 8, -101, 43, 73, -24, -122, 18, 49, -128, -27, 44, 79, 49, -33, -116, 44, 117, -128, -38, 127, -71, 24, 10, 32, -52, -75, 3, 108, 2, -58, 64, -121, 58, 76, -128, 64, 127, -26, -80, -128, -23, 127, 64, -3, -92, 0, 28, -111, -96, 18, 32, 29, -5, 75, 31, -47, 127, 3, -117, 23, -22, 124, 37, -128, 68, 53, 38, 1, -88, -10, 48, 22, -66, 0, 48, 37, -29, -57, -38, 49, 75, -57, 48, 38, -11, 48, -16, -53, -80, 63, 85, -128, 10, -11, -76, 26, 71, -48, -108, 13, 118, 55, -13, 38, -122, -79, 111, 23, -23, 17, 64, -128, 11, 81, -73, -10, -2, -39, -54, 114, -7, -107, 31, 11, 57, 69, 6, -66, 50, 34, -85, -6, -22, -47, 43, 32, 7, -43, -55, 13, 127, 123, -128, -11, 70, -16, -53, -66, -26, 90, -5, -24, 118, -26, -22, -21, 95, -45, -57, 116, 18, -128, -26, 28, -21, 127, 10, -23, -111, -12, 127, -128, -3, 15, 28, 12, 28, -55, -22, -27, 42, 108, -85, -16, -54, 92, 96, -128, -69, 69, 127, 64, -114, -70, -39, 81, 6, 0, 27, -70, -23, 17, -7, -80, 64, -10, -34, 63, -36, -91, 65, -3, -118, 12, 127, -37, -93, 116, 1, -48, 127, -42, -98, 70, 64, -2, -44, -43, 28, 127, 0, -26, 1, -123, -54, 75, 43, 44, -57, -109, 5, 17, 63, 2, 0, 18, -2, 42, 81, -32, -15, 36, -43, 42, -90, -96, 70, 43, -23, 68, 3, 27, 31, -128, -63, 127, 60, -52, 22, -128, 36, 127, -128, -75, 11, 55, 55, -22, -75, 3, 127, 42, -128, -16, 117, -68, 1, 127, -55, -31, 6, 0, -12, -118, 69, 57, -128, 16, 36, 37, 22, -124, 47, 78, -65, -128, 21, 23, 13, 58, -2, -18, -32, 38, 76, 31, -37, -97, 53, -43, -98, 92, -31, 65, 111, -128, -11, 127, -26, -5, 8, -118, -76, 88, -27, 32, 64, -58, 47, -98, -114, 74, 58, -10, -85, 22, 52, 54, 59, -113, 43, 98, -73, 1, -11, -98, 59, -55, -86, 86, -31, -66, 127, 5, -8, -59, -74, 86, 76, -79, 18, -66, 24, 48, -68, 76, 17, -26, -44, -54, 79, -31, -93, 58, 0, -74, -7, 70, 45, 21, 106, -15, -54, 50, 42, -96, 21, -43, -128, 127, 52, -10, 31, -98, -76, 15, -10, 127, -60, -23, 52, 48, -87, -7, 76, -75, 52, 16, -34, 66, 27, -108, -60, 24, -23, -8, 127, -54, -42, 118, 44, -128, -7, 109, -68, -117, -29, 119, 127, -127, -80, 55, 122, -32, -128, 63, 88, 16, 49, -127, -28, 111, -33, -123, -21, 127, 1, -113, 114, 116, -128, 44, -18, -3, 101, -78, 13, 37, -128, 16, 112, -81, -124, 98, 81, -128, -36, 34, 97, -37, -57, 55, -64, -59, 112, 27, 44, -86, -32, 127, 39, -70, -44, 71, -87, -79, 45, -39, -29, 109, -53, -54, 57, 17, -8, 127, 12, -76, 8, -23, 80, 66, -17, -12, -5, -86, -100, 71, 6, 2, 1, -65, -15, -11, 16, 74, 22, 10, 2, -17, -78, 0, -107, 8, -11, -86, 127, 12, -5, -78, 39, 44, 17, 10, -103, 65, -64, -5, 86, -26, -11, -68, 106, 86, -113, -54, 45, -36, -12, 79, -45, 107, 27, -121, 86, 26, -48, -2, 91, -86, -50, 101, -8, -42, -44, 106, -28, -76, 68, 66, 31, 2, -12, -39, -26, -95, 102, -31, -101, 57, 57, 8, -54, 118, 24, 0, -53, 27, -13, -98, -26, 112, 117, -66, -109, -42, 69, 37, -5, 86, 73, 13, -90, -53, 26, -106, 48, 75, -127, 85, 80, -78, -103, 78, 7, -45, 47, -15, -28, -124, 85, 58, -44, 22, -128, 44, 96, -106, -93, -24, 32, 10, 0, 121, 70, -24, 5, -55, -85, 97, -2, -128, 49, 92, -90, -76, 75, 127, 42, -128, 63, 95, -80, 7, -36, -3, 21, -76, -78, 106, 11, -76, -80, 65, 11, 21, 28, -118, -2, 124, 95, -57, -23, -31, -102, 86, 5, -57, 43, -88, -8, 75, -128, -37, 95, 31, -74, -16, -13, 44, 34, 27, -63, -13, 60, -18, -23, 102, -1, -58, 48, -21, -65, 34, 124, -32, -76, 12, -36, -22, 124, -79, -80, 27, 58, 127, 5, -26, -88, 43, -11, -21, 42, -44, -68, 114, 70, -124, 38, -65, 33, 36, -55, -60, 103, 34, -63, -2, 60, 33, -57, -11, -12, -3, -15, -128, 8, 42, -127, -47, 97, 37, 44, 87, -38, -32, 23, -81, -106, 74, 48, -101, -44, 127, -47, 27, 28, -58, 12, -44, 26, -12, -26, 44, 12, -31, 91, 127, -39, -66, 57, 23, -38, -73, -1, -26, -74, 32, 66, -43, -92, -17, 53, 0, -47, 57, -2, 11, -32, 18, 102, -55, -2, -122, 38, -21, -123, 119, -38, 54, 0, 49, 69, -128, 27, 76, -26, 90, -88, -71, 75, -1, 42, -90, 49, -34, 0, 13, 6, -42, -100, 127, 97, -128, 50, 107, -128, -80, 68, 11, 90, 36, -116, 23, 57, 27, 69, -128, 2, 11, -17, 26, 42, -6, -29, 60, -11, -60, 108, -36, -73, -22, 127, -6, -128, 127, 111, -128, -123, 42, 73, 78, 26, -49, -74, -28, 28, 5, 2, 127, -32, -26, -23, 59, -64, -23, 91, -66, 70, -18, -50, -33, -10, 52, -29, -2, 10, -55, 58, 1, -45, -43, -32, 11, 81, 7, -47, -87, 43, 113, -128, -103, 118, 34, -96, 85, -17, 26, 6, -85, 37, 127, -3, -3, -11, 16, -16, -128, 11, 50, 63, -87, 38, 0, -42, 91, 37, -121, 34, 71, -128, -70, 127, 90, -87, 39, -24, -53, 34, -7, -2, 42, -53, -122, 69, 127, -128, -81, 24, 52, 85, 36, -43, -53, -76, -33, 45, 127, -17, -117, 74, 34, -50, 22, -10, 79, 10, -3, -3, 78, -44, 23, 91, -88, 58, -36, -70, -45, 55, 69, -24, -37, -6, -36, 86, 27, -102, -44, 29, 76, -47, 52, 80, -109, -101, -44, 2, 88, 64, -32, -31, 73, -38, 91, -24, -118, 85, 80, -27, -57, 15, 127, 18, -22, -69, -8, 36, 5, 58, 34, -95, -102, 127, -2, -32, 127, -100, -39, 44, -2, 60, -16, -128, 74, 42, -122, -74, 127, 95, -128, -119, 127, -18, -68, 108, -78, 55, 92, -85, -59, -7, 18, -26, -64, -97, -8, 101, -18, 64, 95, -32, -50, -36, -111, 53, 12, -53, 116, -45, -73, 11, 31, 36, 1, 98, 93, -87, -21, 70, -119, -50, 95, -66, -47, 39, 11, 57, 91, -16, -53, 69, -18, 93, -18, -98, 116, 5, 2, 11, -10, 65, -26, -8, 70, -33, -90, 49, -70, -78, 127, -11, 5, 6, -47, 93, -3, -45, -45, 117, 71, -128, -10, 103, -71, -21, 127, -7, -26, -52, 55, -48, -123, 59, 118, 60, -5, -128, -1, -44, -27, 76, -24, -53, 95, 60, 6, -108, 47, 96, -22, -76, 13, -44, -128, 127, 69, -128, 17, 73, -43, 23, 33, -31, 52, -22, -85, 78, 26, -128, 66, -32, -29, 8, -57, 32, 106, -80, -43, 121, 44, -75, -92, 92, 55, -87, 33, -8, -54, 1, 73, 34, -5, -68, -111, 78, 86, -57, -38, -22, 21, -24, -24, -38, 15, -93, -128, 127, 1, -49, 54, 78, 7, -68, -5, -48, -103, 38, 118, -44, 8, 13, -123, 54, -42, -34, 103, -93, -39, 74, 80, -50, -86, 88, 107, -121, 3, 100, 0, -128, -65, 108, -58, -26, 48, 112, 37, -86, -26, 21, 88, -48, -100, 15, 17, 33, 96, 69, -90, 42, -31, -122, 22, 58, 101, -90, -7, 95, -128, 23, 102, -55, -88, 73, 52, -69, 6, -44, 42, 96, -53, -47, -90, 43, 85, -102, -98, 65, 0, 8, 55, -22, 23, 47, -128, -10, 127, -12, -114, -85, 60, -1, 34, 88, 39, -90, -97, 78, 43, 80, -23, -127, 66, 64, 52, -68, 13, -75, 27, -15, -34, 52, -6, -22, -54, 49, 102, -97, -76, 17, -3, 98, -33, 21, 8, -128, 127, 27, -81, -2, -24, 92, -12, 8, -18, -75, -5, 5, 45, -29, 18, -18, 53, -17, -11, -31, 63, 58, -97, -45, 88, 54, -128, -60, 108, 42, -54, 17, 102, -1, -13, -100, -23, 22, -57, -33, 123, 49, -59, -27, 71, -71, -17, 96, -58, -60, 95, -26, 27, -33, -39, 86, 31, -50, -6, -36, -123, -10, 12, -8, 127, 113, -128, -36, 0, -1, 63, -73, -65, 33, 74, 121, -68, -121, 79, 70, -47, -43, 96, -50, -45, 44, -101, 37, 23, -76, 8, 78, 26, -27, 57, 12, -50, 113, 92, -80, -65, 17, 42, -16, 22, -60, -10, -13, 15, 16, 66, 103, -57, -12, -60, -50, 39, 12, 100, 12, -95, 78, 59, -76, -127, -17, 127, -39, -102, 91, 74, -32, -88, 1, -16, 112, 54, -80, 65, 38, -74, -44, 27, -80, -48, 127, -17, -37, -18, -32, 5, 85, -5, 97, -24, -101, 47, 119, -6, -86, 32, -47, -87, 121, 68, -128, 54, -10, 0, 68, 58, -85, -111, 119, 10, -23, 43, 23, 73, -27, -39, 68, -128, 3, 127, -128, -107, 45, 13, 63, 73, -3, -13, -22, -59, -81, 58, -55, -60, 28, 43, -33, -44, 90, -128, 16, 33, -58, 31, -27, -33, 21, 49, 22, -3, 27, 85, 3, 21, 68, 57, -81, -50, 96, -73, -80, 44, -3, 38, 97, -5, -93, -52, 0, 3, 10, -32, 49, 88, -53, -8, 22, -42, -128, -91, 127, 5, -37, -42, 78, 0, 47, -33, -21, 111, -76, -112, 0, 117, 63, -102, -3, 0, 21, 111, -24, -128, -36, 75, -44, 108, 15, 8, 32, -90, -92, 27, 114, -13, -44, -3, 36, -28, -7, 5, -53, -53, 70, 58, 29, -63, 7, -3, -32, 18, -28, -26, 53, 48, -1, 0, -43, 65, -1, -128, 7, 85, 16, -75, -45, 3, 96, 107, -55, -91, -22, 88, -7, -128, 32, 52, -15, -10, 58, 87, -21, -128, -54, 64, 78, 57, 31, -128, 7, 60, -90, -13, -10, 127, 23, -88, -45, 5, 48, 74, 29, -5, -13, -114, 63, -32, -28, 12, -11, 18, -33, -2, 49, 24, 29, -48, -32, 95, -12, 92, 103, -113, -100, -21, 44, 101, 5, -53, 74, 44, -128, -7, 69, 7, 12, -65, -128, 15, 127, -37, 3, -108, 10, 23, -49, 8, -12, 52, 52, -36, -33, 21, 47, -17, -29, -86, -32, 5, 58, 8, -86, -43, 11, 127, 100, -128, -16, -8, 39, 54, -16, 15, -17, -36, 70, -101, 3, 24, -16, 26, 17, -60, -88, 119, -49, -88, 43, 93, 31, 50, 71, -85, -2, -93, -36, 127, -66, -108, 127, 111, -81, -65, 10, -48, -71, 92, 26, 47, 65, -1, -106, -28, -31, 5, 34, -71, 52, 27, 10, -92, -34, 114, 21, -92, 52, -24, -101, 15, 44, 127, -93, 12, 65, -49, -65, 22, 8, -7, 58, -58, 21, 127, 23, -42, -37, -74, 103, -36, -13, 81, -98, -60, 38, 123, -16, -107, -37, 79, 24, -23, 44, -15, -18, -45, 127, 27, -53, -55, 50, 127, -128, -106, 127, 74, -10, -119, 52, 59, -127, 26, -11, -23, 80, -3, -78, -50, -78, 80, -23, -23, 24, 31, 96, -47, -24, 28, 32, -111, 2, 73, -124, 53, 85, -15, -47, -42, -81, 36, 27, -10, 11, 45, -45, -42, 73, 50, 18, -36, -64, 48, -93, -6, 48, 33, -64, -113, 95, 127, -87, -100, 85, 7, -75, 32, 22, 52, 106, -92, -87, -2, 96, 39, 11, -128, -117, 116, 102, 38, -119, -75, 119, -33, 50, -28, -116, 16, 34, 116, -54, 1, -13, 38, 127, -122, -106, 31, 127, -52, -27, 32, -23, 34, 106, -42, -80, 123, 42, -128, 27, 121, -97, -49, -28, -12, 98, -28, -27, -43, -48, 116, 73, -96, -21, 85, -18, -10, 85, -68, -10, 23, -24, 101, 27, -98, -76, 127, -26, -3, -18, 32, 85, -87, -26, -78, -47, 80, 68, 37, -12, 7, -22, -74, 111, 70, -44, 58, 48, -128, -124, 69, 64, -13, -27, -39, 86, 28, -95, 112, -5, -81, 114, 90, -11, -128, 39, 73, -79, -68, -22, 103, 54, -97, 17, -11, -128, 26, 76, -80, 65, 68, -43, -45, -80, 127, 26, -26, -39, -13, 53, -34, 57, -29, -60, 75, 36, -52, -5, 127, -5, -58, 79, -65, -106, 111, 100, -112, -60, 42, 26, -47, 121, 119, -128, 27, 47, -66, -29, 37, -92, -113, 32, 127, -28, -59, 18, 37, 22, -16, -5, 69, -87, -59, 33, 5, -2, 127, 29, -96, -10, 88, 11, -90, 70, 87, -92, -15, 50, 74, -29, -29, 98, -28, -65, -65, 109, 69, -58, -44, -60, -11, 33, 27, 39, 16, 1, 27, -33, 64, 68, -76, -45, 112, -31, -5, 0, -70, -54, 81, -26, -53, 39, -64, -50, 127, -15, 24, 23, -22, -49, -5, -66, -5, 127, -76, 1, -37, 1, -43, -111, 101, 54, -21, 15, -90, 23, 26, 15, 107, -109, 39, 18, -34, -53, 0, 85, -37, 13, -27, -29, 127, 79, -128, -39, 102, 12, -69, -71, 45, 63, -45, -49, -15, 127, 79, -128, -42, 127, 34, -128, -86, 109, 60, -6, 23, -116, -57, 127, 13, -117, -23, 39, -3, 24, 114, 66, -128, -70, 24, 85, 108, -73, 2, 80, -121, -29, -24, 33, 54, 21, 33, -60, -47, -16, -15, -11, 43, 60, -48, 90, 79, -103, -68, 108, 55, 13, -23, -29, -87, 32, 22, 29, 116, -128, -2, 26, -24, 87, 29, -128, -6, 96, -29, 59, 24, -57, -128, -44, 33, 0, 127, 63, -116, -87, 33, 127, 43, -21, -88, 8, -18, -33, 28, -59, 12, -26, -1, -22, -74, 58, 5, 52, -63, 26, 80, -5, -63, -15, -80, -16, 127, -121, -69, 55, -28, 101, -21, 66, 48, -78, 64, -107, -58, 106, 29, -76, -55, 59, 74, -16, 68, 69, -128, 55, 65, -48, 39, -128, -12, -29, 47, 74, -119, -53, 127, -11, -5, 111, -123, -71, 85, -47, -1, 127, 3, -1, 27, -60, -118, -10, -27, -17, 69, 6, -12, 127, 114, -128, -102, 127, -23, 79, -10, -91, -3, 127, 31, -39, 52, -38, -123, -18, 111, 10, -79, 0, 63, -39, 114, 58, -103, 54, 8, -43, -128, 47, 92, -128, 73, 106, -75, -128, 49, 112, -106, 13, 53, -18, -34, -28, -28, 17, 65, 49, -128, 36, 17, -73, -11, -1, 15, 80, 0, 55, 6, -103, 93, -57, -60, 116, 55, -1, -43, -70, -5, -95, -23, 57, 60, 53, -2, -128, -42, 114, -85, -11, 100, -53, 49, 33, -66, -112, -17, 127, -107, 17, 17, -1, 96, -74, -63, 36, -23, -74, -1, -18, 6, 90, 5, -108, 27, 33, -52, -44, -7, 60, 78, -128, 59, 97, -59, -37, 16, -91, -39, 127, -124, 7, 119, -128, -12, 65, 71, -91, 22, 38, -79, 18, -6, -43, 91, 127, -39, -128, -44, 127, 55, -128, 73, 85, -55, 1, -88, -6, 90, 5, -74, -128, 66, 53, -116, 1, 127, 93, -121, -22, -2, 17, -54, 0, 111, 3, -42, -66, 60, 48, -116, -16, 81, -73, -68, 78, -59, 39, 37, -108, 78, 127, -121, -50, 59, -36, 86, -6, -79, 127, 85, -116, -15, 59, 39, -106, -49, 28, 26, -18, -55, -34, -5, 34, 66, 38, 59, -2, -116, 127, 23, -68, 74, -43, -128, -21, 117, 68, -80, 26, 33, 54, -100, -118, 127, 118, -87, -101, 32, -27, 55, 91, -117, 17, 95, -58, -117, 18, 127, -98, -45, 22, 52, -23, -8, 55, -76, -70, -8, 59, -75, -111, 127, 1, -93, 96, -15, 17, 111, -33, -17, -8, -79, 81, -21, -121, 53, 37, 34, -29, -6, -39, 23, 12, -32, 2, -64, -57, -34, -42, 11, 65, -16, -58, 98, 24, -13, 71, -128, -17, 68, 45, -80, 18, 98, -71, -111, 16, -2, 106, 102, -39, -114, 10, 23, -116, 45, -29, 23, -39, -42, 3, 33, 75, -87, -44, -12, -48, 37, 29, 45, 74, -121, 15, 64, 7, -87, -13, -3, -55, 78, -37, -47, -2, 3, -11, 78, 0, -11, 70, -10, -87, 108, -6, 18, -10, -18, -23, -27, -12, 37, 6, -95, 127, -27, 0, 116, -81, -23, -45, 76, 2, -52, 0, 8, 87, -44, -90, -48, 127, 96, -92, -123, 66, 100, 32, -128, -34, 39, 7, 64, 27, -15, -38, -32, 6, -49, -53, -23, -64, 98, 1, -29, 12, 32, -31, -54, 127, -5, -128, 127, 121, -92, -24, 10, -108, 38, 47, -6, -117, -58, 111, -57, -43, 79, 107, -88, 60, 21, -79, -33, 127, 57, -96, -32, -44, 70, 24, 90, 32, -121, 39, 17, 5, -13, -106, -48, 54, -26, -44, 117, 28, 11, 26, -23, -86, -1, 86, 91, -32, -24, 45, -79, -81, -16, 64, -11, 21, -87, -36, 87, -8, -26, -29, 27, 127, -21, -52, -6, -15, 57, -111, 65, 37, -52, 8, -34, 80, 64, -122, -65, 92, -44, -116, 18, 114, 63, -22, -60, 28, -69, -112, 50, 79, -26, 47, 16, 3, -34, 39, -22, -128, 127, -7, -63, 65, 11, 55, -50, -36, -32, 79, 1, -66, 101, -7, -128, 49, 0, 5, 27, -58, 29, 45, -128, -111, 127, 36, 28, -108, -36, 38, -43, 59, 39, 28, 73, 42, -91, -92, 34, 74, -63, 69, -3, -97, 93, 43, 68, 60, -128, -17, 54, -65, 37, 75, -39, -32, 0, 18, 34, 75, 6, -36, 107, 15, -17, 3, -54, -78, 90, 96, -55, 13, -31, -28, 53, 7, 3, -54, -43, -70, -64, 127, -22, -55, 66, -31, 44, 12, -42, 70, -108, 16, 1, 28, 1, 12, 1, -42, 92, -107, -59, 66, 86, 21, 6, -34, -85, 63, -80, 48, 107, -128, 38, 116, -75, -93, -29, 0, 98, 63, -128, 39, 47, -114, 38, 80, -112, -93, 70, 127, -86, -21, 26, 52, -10, -101, 47, 81, 76, -65, -45, 48, -23, -36, 28, -68, 47, 113, -101, -31, 38, -28, -21, -68, 74, -12, -128, 127, 6, -103, 121, -47, 29, -49, -109, 50, 24, 52, 103, -95, 37, 26, -13, -15, 21, -15, -53, 57, -59, 64, -3, -128, 66, 127, -90, -55, 0, -11, 52, 17, 38, -45, 23, 38, -86, 49, 38, -69, -74, 6, 53, -66, -101, 70, 93, 33, 22, -128, -22, 13, -60, 127, -24, -26, 101, -63, -95, -53, 123, 71, -64, -13, -90, 10, 34, 23, 29, -59, -13, 127, 60, 7, -128, 11, 48, -6, 34, -85, 73, -37, -58, 127, -108, -32, 109, 24, -128, 44, -36, -128, 127, 73, -38, 28, -114, 47, 21, -71, 123, -23, -117, 69, 13, -49, 29, 73, 75, 12, -18, -47, 27, -90, -36, 118, 11, -127, 28, -60, -69, 127, -65, -118, 107, 92, 24, -37, -57, 78, 45, -128, -80, 127, 50, -98, -101, -32, 7, 127, 96, -43, -70, -12, 86, -128, -29, 127, -65, -52, 76, 21, -106, 43, 38, -28, -39, -49, -34, 100, -2, -127, -1, 114, -28, -87, 47, 47, -5, 23, 2, 121, 117, -100, -69, 65, -17, -128, 38, 114, -49, -79, 0, 64, -66, -96, 66, 68, -8, -128, 52, 17, -96, -1, 127, 10, -121, -6, 90, 8, -33, 80, -47, -31, 13, 80, -17, 5, 107, -128, 5, 88, -57, -24, -1, 71, 12, -128, 26, 33, -103, 26, 65, -63, -6, 31, -128, -74, 34, 100, 48, -29, -15, 32, 71, -32, -63, -59, 24, 53, -38, 0, -11, 100, 88, -47, -3, -11, -128, 52, 32, -33, 48, -36, -45, 73, 5, -34, 114, -10, 52, -34, 8, 3, 28, 50, 2, -65, 22, -2, 0, 118, -54, -23, 39, -80, -17, 47, 81, -33, 48, 86, -79, -78, -87, 71, 109, -128, 23, 23, -92, 45, -1, 53, 17, -128, -6, 53, -37, 127, 0, -47, 49, -3, -81, -64, 113, 11, -48, -1, 29, -8, -50, 2, -79, 59, 23, 38, 85, -128, -50, 23, 71, 81, -119, -42, 127, -10, -18, -86, 2, 10, 65, 0, 16, 118, -96, -45, 15, -93, -16, 57, 73, 44, 8, -15, -70, -81, 74, 23, -54, 127, -3, 6, 21, -70, -45, 15, -50, 112, 45, -79, -54, -23, 118, 98, -103, -93, 81, 90, -70, 12, 117, -6, -118, 10, 6, -10, 43, 28, -17, -22, -8, -128, 36, 21, -7, -59, 48, 74, 17, -81, -119, -3, 69, 114, 42, -65, 10, -52, -91, -27, 127, -24, -5, 8, 15, -28, 28, 48, -128, 63, 34, 31, 60, -127, -59, 85, -8, 102, 127, -128, -96, 39, 5, 90, 102, 36, -128, 0, 15, -65, 107, -43, -38, 69, -2, -54, 70, -3, 3, 71, 5, 28, -73, -68, 102, -18, -34, 81, -96, -22, -52, -12, 127, -76, -101, 121, -8, -54, 68, 16, 34, -44, 3, 127, -27, -8, -101, -69, 15, 79, 117, -7, -66, -70, -23, 45, 86, 74, -90, 42, 18, -111, 17, -3, 8, 52, -102, 31, 127, -66, -128, 32, 87, 10, -33, -54, 32, 43, -10, 17, -52, -8, 39, 57, 32, -33, 71, 108, -128, -128, 127, 58, -107, -16, 87, 58, -128, -128, 127, -17, -18, 127, -16, -112, 2, 127, -52, 5, -7, -11, -5, -50, 114, -15, -3, -50, 0, 57, -98, 59, 60, -116, -13, 127, 2, -128, 75, 37, -122, 0, 50, 12, -70, -101, 101, 68, -128, -65, 106, 15, 36, 45, -45, -26, -86, -17, 100, 49, -128, -114, 127, 78, -93, -70, 96, 109, -60, -24, 10, 33, -57, -71, 79, 48, -37, -15, -17, 5, 52, -113, -93, 121, 111, -3, -103, -90, 28, 26, -28, 45, 27, 81, -73, -33, 127, -7, -103, -28, -3, 107, -45, -29, 1, 65, -11, -5, 16, 0, -10, -87, 86, 8, 2, 17, -108, -48, -58, 98, 92, -121, -53, 127, 98, -128, -60, 109, 29, -28, -118, -88, 108, 11, -2, 78, -100, -128, 103, 95, 3, -107, -107, 123, 103, -128, 5, 26, -6, 59, 93, -113, -6, 7, 68, 58, -119, -2, 33, -36, -21, 93, 8, -113, -7, 36, 127, 5, -124, 69, -12, -88, 127, -5, 2, 45, -88, -21, 81, 38, 6, -21, -18, -29, 16, 15, 38, 53, -128, -39, 47, -7, 0, 68, 13, -60, 96, -38, -2, -37, -128, 127, -10, -16, -23, 43, -2, -80, -8, 91, 93, -32, -109, -39, -10, -59, 6, 59, 3, 0, 127, 0, -17, -43, -65, 127, 8, -1, -22, -108, -8, 47, 18, 8, -1, 27, 22, 5, 80, -17, -79, 59, -18, 7, -32, -18, 85, -78, 7, 57, -90, -34, -54, -76, 98, 12, -80, -3, 42, 71, 1, -17, 90, -8, -17, -90, -97, 34, 95, 100, -12, -128, 44, -2, 43, -38, 6, 97, -88, 5, 17, -124, 1, -26, -3, 48, -1, 49, -7, 29, -74, 44, 1, -122, 88, -5, -33, 106, -1, -118, 90, 12, -81, 81, 42, -70, 74, 17, 55, -23, -112, 107, 27, 5, 27, 12, -123, -88, 96, 65, -111, 50, 79, -97, 86, -49, -50, 18, 64, 80, -128, -22, -38, 7, 7, 11, 71, 28, 21, -69, 36, 66, -128, -48, 103, 64, -88, 10, -53, 38, 45, -128, 58, 127, -73, -52, -48, 71, 103, -128, 38, 6, -28, 114, -36, -29, -49, -79, 50, -16, 48, 34, 58, 22, -43, -15, -47, 88, -55, -70, 96, 0, -47, -42, 22, -68, -85, 127, 118, -32, -43, -17, -128, -18, 106, 17, -81, -101, 127, 85, -128, -11, 127, 42, -17, -70, -88, -12, 27, 32, 49, -74, -80, 34, 80, -112, -22, 127, 6, -80, -15, 15, -91, 38, -33, -121, 91, 59, -87, 29, 7, -38, 127, 108, -7, -60, -76, -43, -45, -17, 21, 13, 85, 53, 17, -32, -3, -12, -36, 33, 102, -85, -85, 63, -32, 57, 57, 5, 87, -38, -128, -38, 118, 108, 34, -66, -70, -8, 66, -1, -59, -109, 65, -7, -23, 52, -8, -58, 48, 91, -54, -26, -128, 78, -12, -128, 107, 54, 27, -24, 47, 22, -97, -10, 13, -7, -66, 122, 117, -128, 5, 88, -109, 18, 91, 23, -124, -33, -3, 123, 3, -28, 65, -95, 17, 60, -70, -73, -16, 127, 36, -128, 43, 127, -44, -128, -3, 107, -47, -43, 108, 71, -7, -11, -86, -32, 42, -32, 48, 6, -87, -63, 29, -10, 39, -3, 60, 107, -128, 32, 63, -39, -128, -28, 127, -13, -32, -73, -43, 117, -2, 32, 10, -128, 50, 103, -23, -103, -43, 54, 80, -13, -37, -88, 26, -27, -59, 76, -79, 28, 78, -128, 18, 109, -45, -48, -18, -47, 53, 50, 36, -127, -29, 79, -53, -8, 26, 119, 1, -47, -1, -31, -10, -28, 79, -36, -26, 8, -96, -53, 49, 127, -70, -128, 127, 81, -42, -106, 87, -18, -21, 93, -116, -60, 13, 27, 43, 10, -28, -68, 15, -21, 75, 121, -80, -18, -31, -55, 0, 48, 3, 16, 11, -34, 44, -50, -66, 32, 42, -32, 44, 10, -75, -37, 127, 53, -42, -6, -48, -38, 101, 80, -92, 1, 65, 44, -71, 64, -42, -39, 85, -6, -33, -59, 127, 124, -128, -88, 22, 98, 12, -128, -26, 127, -53, 68, -7, -44, 29, -47, 50, 79, 2, -52, -96, -44, 23, 29, -32, -7, 127, -1, -26, -107, -8, 119, -117, -101, 38, 85, 112, 1, -55, -93, 1, 108, -74, 23, 31, -32, 113, 50, -128, 0, 28, -27, -74, -81, 33, 69, 44, -36, -47, 49, 33, 78, -49, -49, 113, -60, 22, 47, -128, -2, 127, -37, -114, 109, -44, -50, 64, -66, 28, 112, 69, -128, -29, 24, -42, 119, 42, -7, -116, 48, 8, -49, 96, -28, 54, -8, -38, 66, -118, 3, 33, -122, -1, 117, -64, -15, 33, 10, 52, 32, -53, -12, 93, 29, -39, 38, -27, -113, 63, 32, 49, 21, -26, -29, -123, 79, -29, 34, 96, -118, 29, -24, -39, 127, 37, -117, -70, 103, 29, -49, -59, 28, -74, -103, 91, 60, 49, 10, -59, -63, -70, 42, -10, -66, 21, 43, 127, -38, -97, 90, 38, 47, 10, -10, 12, -64, -75, -26, 49, 127, 37, -42, -15, -128, -95, 85, 111, -74, -38, 80, 37, 23, -96, 58, 93, -128, 93, 23, -116, -34, 124, 59, -17, -42, -65, 24, 69, -24, -31, -55, -7, 57, -68, -13, 85, -47, 37, -2, -70, -32, 88, 102, -60, -16, -13, -103, 74, 24, -48, -70, 18, 44, 21, -29, 33, -53, -128, 127, 97, -36, -119, -26, 50, -8, 93, -81, -5, 101, -54, -109, 100, 1, 23, 27, -128, 39, 101, 57, -128, -60, 16, 65, 98, 7, -128, 16, -12, -85, 101, 92, 12, -48, -113, -47, -6, -7, 45, 101, 39, -38, -17, -36, -128, 57, 0, -107, 45, 127, -78, -53, 38, -28, 1, 2, 10, 57, -31, 5, 109, 36, -78, 8, 17, 6, -91, 22, 127, -74, -53, 59, -63, -42, 32, -16, -36, 44, 32, -128, 63, -12, -44, 50, -31, 92, 1, -32, -48, 0, 109, 28, -128, -85, 69, 78, -128, 10, 91, -128, -12, 45, 109, 37, -26, -33, -93, -10, 39, -48, 0, 52, -31, -76, 114, 70, -13, -60, -75, -32, 127, 1, -128, 28, 96, 66, -111, 17, 45, -8, 24, 1, -128, 17, 71, 31, -66, 8, -10, 3, -70, 17, 24, -70, -68, 3, 31, 93, 57, -75, -117, 58, 124, -121, -109, 85, 127, -85, -95, 54, 127, -100, -100, 127, 33, -58, 37, -128, 1, 58, -128, 127, 24, -74, 27, -31, 64, 27, -116, 6, -15, -34, 34, -47, 42, 42, 5, -10, -8, 47, 11, -80, 0, -98, -32, 87, -128, 15, 117, 10, -128, 34, 111, -87, -48, -16, 101, -13, -124, 36, 2, 34, 117, -11, -21, -17, -85, 13, 127, 39, -128, 43, 10, -103, -22, -10, 127, -34, -24, 78, 6, -12, -81, 2, -68, 45, 121, -128, -85, 26, 47, 33, 31, -33, 73, -21, -42, 127, -36, -73, 29, 45, -59, -93, -24, 93, 29, -85, 91, 127, -36, -79, 12, -66, -66, 127, -52, -80, 7, 39, 58, 3, 43, 58, -39, -58, -75, -29, 74, 64, 31, -92, -2, 1, -7, 86, 43, -7, -8, -43, 16, -12, 73, -21, -49, -2, -33, 95, 28, -57, -63, 121, 80, -49, 2, -74, -79, 106, 8, -34, -7, -95, 70, 102, -123, -114, 50, 118, 11, -128, -39, 59, 27, -17, 49, 113, -74, 3, 8, 6, -86, -21, 97, 26, -81, -34, -15, 36, 15, 23, -28, 38, -80, -93, 127, -27, -73, 26, -23, -28, 48, 48, -18, 44, 18, -128, 43, -22, 53, 1, 15, -60, 11, 80, -3, -79, -90, 10, 127, 42, 2, -73, -32, -45, 29, 87, -42, -52, -42, 127, 31, -24, -17, 63, 8, -128, 127, 1, -128, 127, 12, 3, 64, -128, -27, 92, -53, -2, 70, -98, -75, 108, 5, 3, 29, -128, -22, 17, -15, 48, 97, 5, -128, -34, 101, 33, -54, 15, 66, -44, -22, -33, 10, 50, -6, 118, -74, -8, 85, 6, 27, -23, -63, -79, 31, -22, -21, -43, 26, -69, 36, 93, -52, 17, 26, -128, -60, 2, 86, -47, -11, 31, -69, 127, 29, -88, 54, 7, -108, 2, 66, -48, 10, 13, 68, -7, 23, 15, -21, 18, -22, 5, -21, -22, 55, 13, 24, 109, -12, -87, 93, 111, -107, 11, 45, -21, -87, -32, 16, -16, 86, 32, -75, -102, 101, -37, -79, 93, -11, 54, -107, 16, 28, -118, 127, 32, -114, -18, 6, 70, 7, 68, -16, -45, 70, -107, -15, -3, 36, 117, -53, -54, 33, -98, 39, 81, -106, -49, 17, 102, -47, -55, 90, -6, -16, 21, -111, 66, 117, -128, -37, 8, -32, 121, 78, -13, 3, -116, -128, 95, 10, 8, -11, 54, 68, -128, 22, -3, -22, -8, 108, 64, -97, 18, -57, -63, 50, 8, 127, -49, -71, 66, -29, 50, -7, -66, 88, 5, -2, 68, 48, -2, -100, -78, 106, -18, -50, 75, -13, 60, 34, -85, -7, 127, 49, -97, -106, -32, 127, -18, -52, 28, 58, 50, 27, 17, -23, -81, 75, -59, 16, 93, -31, -113, 45, 39, -102, -34, 127, 17, -3, -32, -12, -23, -32, 68, 55, -23, 3, -8, -11, 87, -31, 34, -37, -119, 86, 114, -65, -55, 107, -58, -98, 107, 5, 63, 95, -107, -128, 90, 111, -18, -128, -37, 127, -60, 0, 11, -33, -27, 33, -55, -75, 32, 127, 0, -117, 65, -21, 13, 123, 31, -74, 13, -59, -16, 66, -100, -93, 116, -42, -118, 127, -6, -21, 60, -15, -32, -59, -17, 116, 90, -128, 27, -54, -87, 58, 3, 93, -12, 8, 38, -97, -12, 64, 42, -60, -2, -26, 42, 58, -58, 79, -32, -13, 27, 59, -60, 24, -31, -49, 112, 68, -21, -58, -123, 90, 114, -128, 5, -12, -87, 54, 65, 12, 69, 76, -58, -112, -64, 13, 127, -8, 42, 59, -32, -108, -13, 122, -128, -13, 39, 8, 42, -117, -17, 117, -58, -58, 127, 59, -128, 47, 86, -70, -116, 38, 36, 2, 42, -57, -128, 32, 127, 17, -106, -16, -34, -88, 114, 8, 11, 103, 7, -122, -128, 21, 127, -73, -69, 127, 17, -38, -8, -8, -78, 73, -21, -8, 65, -116, -36, 85, 53, -106, -8, 0, -113, 127, 27, -29, -34, -73, 124, -16, -17, 111, -28, -44, 66, 57, -102, -27, 49, 65, 75, -59, -36, -59, -16, 37, 1, 79, -74, -58, 5, 92, 55, -128, 45, -49, 28, 123, -128, -43, 127, -16, -128, -26, 127, 48, -21, 24, -128, -87, 122, 97, -10, -114, -78, 1, 102, 58, -116, -88, 29, 68, 119, 34, -80, -32, 36, -60, -44, -65, -74, 101, 95, -92, 43, 32, 7, 10, -98, 50, 60, -128, 32, 80, -91, -76, -50, 43, 127, -52, -74, -7, 68, 32, -109, 38, 31, -60, 127, 101, -128, -97, 66, 127, -53, -88, 52, -13, 102, 91, -128, 27, 127, -128, -26, 76, -59, 34, 90, -98, 34, -16, -75, 71, 26, -28, -108, 90, 64, -128, 53, 106, -113, -75, 103, 29, -48, 103, 5, -124, 57, 63, -128, 37, 101, -17, -103, 93, -12, 13, -15, -113, 28, 85, 73, 23, -128, 17, 80, -45, -128, 0, 90, -76, 59, -26, -13, 127, 44, -128, -92, 127, 52, -85, -23, 17, 96, 5, -86, -32, 52, 75, -31, 49, -15, -71, 107, 37, -85, 50, 22, -49, 127, 58, -128, 29, 63, 1, -21, -26, 12, 22, -88, -68, 127, 1, -79, 33, 37, -28, -29, -86, -66, -29, 127, 29, -128, 49, 101, -85, 49, 93, -128, 39, 15, -60, 17, 112, -92, 28, 53, -45, 18, -2, -124, 22, 28, -5, 24, -66, 15, 5, 24, 64, -55, -29, 127, -55, -10, 29, -88, 28, -32, -10, 17, -6, 60, 5, -93, 21, 23, -128, 27, 55, 0, 38, -119, -86, 64, 81, -37, 28, 55, -22, -81, -116, 0, 53, 24, -43, -49, -7, -3, 93, 93, -15, -91, 38, 18, 12, 29, -111, 57, 6, -22, 47, -91, -112, 127, 90, -59, -74, 3, 47, -66, -68, 111, 45, -44, -42, -112, -64, 127, 0, -2, 21, 12, 60, -128, -79, 108, 70, -53, -31, -36, -26, 26, 49, -1, -31, 23, -29, 92, -22, 48, -6, -59, 127, 70, -116, -50, -8, 17, 22, 18, -15, 74, 2, 57, 73, -108, -11, 8, 55, -96, 2, 0, -36, 21, 7, 66, -5, -32, -38, 23, -15, -13, -45, -26, 87, 15, 36, 23, 2, 28, 12, -22, -93, 69, 23, -128, 13, 22, 52, 18, -39, 23, 28, 57, 13, -128, 8, 39, 24, -60, -70, 38, 100, -2, -37, 127, -17, -11, -17, 36, 5, -128, 45, 112, -101, -86, 127, 28, -93, 7, 79, 0, 0, -66, -54, 45, -7, -76, -48, 45, 37, -3, 32, 108, -38, -15, 64, -5, -58, 76, 0, -21, -71, -90, 121, 5, -38, 54, 65, 1, 32, -29, -112, 64, 78, -29, -86, -44, -76, 42, 117, -92, 27, -47, 47, 124, -96, -64, -16, 63, -16, -128, 71, 88, -107, -24, 124, -8, 0, -6, 43, 0, -7, -76, -69, 122, -75, -124, 88, 22, 52, -12, -15, 49, -29, 18, 16, 70, 69, -29, -42, -81, 34, -21, 13, 64, -76, -36, -59, -26, -12, -3, 127, -73, -49, 70, 58, 6, -86, -49, 81, -63, -32, 33, -2, 70, 2, 3, -33, -39, 24, -65, 74, 8, -54, 79, -59, -80, 52, 55, 6, -11, 39, -18, -33, -39, 81, -5, -1, -33, -23, 48, -65, -66, -71, 127, -47, -36, 124, -50, -88, -5, 102, -64, 33, 13, 24, 109, -98, -98, 29, 107, 24, -128, -27, 22, 28, 1, 48, -3, -1, 13, -91, -36, 124, -26, -106, 127, -73, -116, 108, 13, 12, -7, 1, 16, 15, 127, 74, -92, -113, -8, 44, 91, -22, -13, -63, -108, 37, -2, 87, -13, 21, 127, -81, -31, -28, 31, 44, -93, 50, 101, -90, -112, -42, 111, 18, -55, 97, -39, 48, 98, -81, -85, 74, -52, -66, 22, 16, 86, -32, 73, 38, -22, 6, 8, -64, -128, 93, -8, -53, 93, 102, -7, -49, -117, -32, 127, -59, 31, -49, -128, 127, 44, -74, 17, 23, -6, -8, 29, -119, 7, 71, -48, -23, -55, 11, -78, -15, 54, -76, 86, -49, -90, 109, 78, -92, 43, 48, -101, 44, 7, -70, 10, -59, -95, 60, -27, 96, 18, -128, 27, 38, 117, 95, -15, -118, -6, -42, -102, 57, 57, 97, -42, -42, 27, -101, 85, 18, -18, -26, -69, 39, -66, -27, -8, 15, 127, -68, -65, 32, -2, 76, 18, 102, -3, -111, 36, 0, 23, 48, 5, 70, -52, 13, 17, -128, -33, 113, 58, -86, -49, 21, 127, -1, -57, 91, 2, -108, 53, 73, -127, 38, -47, -53, 112, -39, -6, -69, 8, -13, 8, 3, -78, 8, 28, 117, -34, -33, 31, 54, 13, -48, -100, 11, 127, -22, -95, 13, 88, -71, -45, 12, -18, 81, 95, -107, -71, 118, 0, 52, 71, -128, -57, 24, 18, 87, 91, -47, 38, -53, -107, 87, 73, -70, -100, 86, 103, -57, -97, 54, 68, -28, 15, 37, -123, -24, 127, -59, -103, 13, 43, -21, 23, 100, -48, 11, 127, 8, -43, 17, -128, -98, 116, 92, -53, -12, 0, -65, -39, 79, 106, -2, -127, 5, 66, -50, -49, 38, 87, -39, 1, 100, -93, 15, 1, -90, 17, 21, -27, 3, 49, -8, 21, 127, -116, 17, 90, -85, -76, 79, -34, 57, 45, -128, 53, -44, 15, 118, -34, -73, -36, 16, 34, 47, 127, -13, -52, -31, 36, 54, -55, -91, -69, 16, 53, -7, 127, 92, -103, -103, 34, 79, -75, -74, 127, 92, -128, -12, 74, 10, 27, -12, -2, 31, 22, -31, -98, 0, 127, -92, -79, 109, -3, -33, 73, 17, -52, 47, -24, 42, 58, -21, -75, 13, 58, -128, -27, 107, -23, 15, -59, -113, 32, 116, 54, -128, -29, -10, 54, 52, -93, 112, 111, -109, -101, 48, 108, -16, -122, 127, -5, -29, 80, -50, -26, -15, 42, -86, -44, 69, -58, 71, 71, -57, 10, -7, -2, 95, -50, -124, 11, 52, 123, -97, -3, -7, -16, 71, -13, 15, -11, 29, -23, -66, 10, 127, 52, -128, -73, 38, 101, -17, 80, -23, -23, 59, -1, -36, 0, 127, -47, -18, 18, -58, 79, 127, -100, -114, 68, 81, 16, 23, -86, 23, 92, -106, -24, 8, -52, 15, 16, -128, 49, 68, -128, -5, 127, -7, -73, -37, 0, 76, 55, -31, 6, -39, -34, 107, -38, 0, 10, -128, 54, 124, -128, 11, 50, 28, -8, -128, 97, 17, -88, 96, 97, -95, 58, 36, -50, -44, 8, 85, 0, -113, -60, 38, 23, 37, -52, -128, 70, 127, -128, -70, 127, -55, -91, 21, 127, 13, -128, 71, 65, -76, -29, 26, 45, -22, 95, -34, -36, 93, -87, -3, 127, -32, 2, 3, -111, -16, 71, -70, -36, 127, -6, -128, 114, 36, -128, 88, 85, -128, -37, 12, -7, 45, 7, -128, -91, 127, 2, 6, 8, -52, 127, -49, -33, 127, -13, -128, -22, 91, -47, 75, 8, -22, 102, -73, -100, 15, 44, -3, 64, 122, -22, -121, 53, 15, -80, 76, 98, -91, -92, -26, 75, 13, -45, 31, -10, 127, -6, -64, 27, -2, -17, 48, 127, -128, 26, 0, -87, 39, 3, 113, 112, -49, -16, -11, -128, -47, 97, -37, 38, 119, -97, -81, 127, -7, -80, -21, -6, 109, 28, -29, 73, 0, -128, 68, 81, -128, 78, 127, -128, -95, 127, -33, 53, 58, -34, 39, -17, -128, 53, 10, -128, -10, 127, -37, 10, 12, -49, 127, 69, -29, -69, 27, 0, -31, 65, -73, 1, 92, 68, -38, -33, 0, -21, 8, -75, -5, 59, 80, -6, -81, -43, 36, 39, -128, 49, 18, -113, 127, 108, -52, -70, -75, 6, 106, 5, 21, 0, -2, -64, -45, 8, -65, -13, -1, 121, 22, -37, 3, -8, -15, 98, 60, -8, -57, -21, 8, -27, 22, -50, -33, 0, 53, 1, -22, -16, -107, 49, 12, -76, -2, 127, 45, -100, -68, 96, -10, -12, 24, 2, 112, -21, -74, 58, 0, 64, -13, 42, 5, 38, -39, 1, 29, -122, 55, 16, 36, 65, 15, 17, -42, 2, -12, -111, -65, 96, 100, -109, -116, 127, 31, -33, -60, 7, -6, -29, 42, -10, 127, 15, -128, -8, 49, 58, -16, 54, 45, 7, -54, -52, 58, 98, -79, -88, 17, 29, 127, -100, -24, -2, 88, -24, -6, -3, -6, 122, -87, 23, -66, -54, 71, -36, 49, 69, -8, 22, -52, -78, 63, 68, -15, 92, -29, -43, -27, -1, 127, -103, -48, 87, -75, 7, 70, 52, -27, -113, 37, 103, -128, 2, 15, -55, 102, 33, -128, -21, 90, -38, 13, 100, -2, -11, -5, 16, -88, -2, 5, -79, -53, -32, 127, -13, -55, 76, -76, -53, 127, 96, -128, -112, 127, 43, -32, 33, -55, 0, 127, -17, -49, -34, -32, 0, -15, -6, 26, 93, -63, 64, -17, -107, 127, 113, -128, -66, 54, -11, 12, 0, -50, 63, 2, 48, -91, 22, 50, -116, 11, 22, 85, -90, 16, 18, -58, -29, 22, 103, 10, -49, -29, 23, 0, -63, 1, 64, 3, -128, -60, 49, 36, 22, -86, -73, 102, 21, -80, -1, 106, 44, -10, -8, 7, -22, 42, -81, -22, 33, 52, -21, -128, 73, 12, 47, -39, 45, 80, -5, -103, -117, 75, 112, 21, -39, -128, 7, 11, -44, 121, 64, -8, -66, -58, 29, 108, -68, -21, 53, -2, 0, 43, 1, -127, -57, 79, 10, 124, -37, -109, 50, 22, 103, -34, -69, 93, 1, 52, 53, -52, -2, -15, 127, 44, -107, -11, 15, 21, 80, 38, -128, -32, 114, 18, -43, 3, 66, -43, -47, -106, 45, 118, -113, -48, 114, -47, -6, 86, -3, -128, -85, 22, 52, 0, 78, 80, -63, 85, -74, -97, 127, -54, 5, 50, 15, -47, -78, 116, 87, -12, -18, -43, -29, 64, 43, -114, -98, 90, -17, 74, 73, -128, -101, 127, 1, -53, 38, -7, 0, -23, 50, -63, -27, 24, 18, -42, -10, 74, 39, -101, -50, 50, 31, 52, -81, -38, -28, 16, -2, -16, 59, 80, -15, -70, 39, 37, -128, -54, 60, 39, 55, -86, -128, 58, 117, -1, -12, -70, -42, 57, 3, 42, -90, -76, 127, 3, 16, -101, -93, 44, 57, 81, 74, 31, -128, 0, 102, -103, -87, 27, -8, -17, 119, -31, 8, 38, 16, -34, 0, -33, -114, 54, 17, -26, 114, -73, 28, 98, -128, 73, 93, -117, -21, 52, -53, 10, 21, -87, -60, 113, 55, -102, -85, 38, 64, 59, -119, -31, 54, 57, 48, -91, -63, -68, 101, -2, -111, 100, 108, -119, -23, 64, -16, -75, -17, -17, -33, 11, 70, 38, -71, -7, 127, -42, 0, 23, -117, 100, -59, -28, 127, 17, -128, -71, 2, -17, 101, 6, 49, 8, -59, 13, -59, -26, -50, 97, 69, -117, -66, 3, 122, -24, -34, 58, -13, -45, -73, 88, 1, -103, 47, -6, -52, 93, 33, -80, -102, 0, 127, -81, -127, 116, 111, -50, -109, -55, 76, 127, -58, -21, -33, -50, -13, 127, -44, 0, 49, -87, 78, -106, 28, 73, -80, -32, 31, -15, 60, 44, -47, 7, -6, -15, -73, -11, -34, -5, 66, -128, 16, 38, 18, -69, -2, 127, 5, -57, -34, -57, -92, 52, 34, -95, -7, -13, 48, 127, -60, -65, 66, -55, -24, 70, 106, 34, -128, -45, 80, -60, -5, 47, 6, -15, 7, -3, -10, 44, 127, -100, 17, 11, -13, 22, -49, -54, 16, 127, 29, -53, -109, -36, 88, -18, 2, 13, -100, -85, 0, -6, 29, 109, -11, 6, 60, -33, -7, -128, -103, 127, -28, -116, 33, -11, 85, 100, -98, -74, 118, -34, 69, -42, -39, 127, -31, -47, 5, -100, 44, 121, -128, -101, 93, 69, -127, 17, 87, -123, 69, 119, -128, -73, 32, 48, 27, 87, -48, -37, 127, 16, -86, 16, 26, -128, 7, 27, 11, -37, -39, 47, -53, -127, -23, 48, 122, -33, 37, 8, -107, 96, -27, -69, 127, -45, -31, -10, -96, 118, 85, -128, 21, 50, -100, 57, 92, 43, -112, -10, 34, 45, -13, -6, 55, -70, -128, 42, 114, -128, -85, 38, 127, 2, -60, 85, 7, -103, -86, 127, -36, 8, 119, -47, -128, 71, -18, -12, 85, -100, -32, -13, -22, 127, -53, -101, 109, -11, 75, 3, -111, 127, 12, -128, 16, -16, 127, -26, -90, 22, 116, 7, 0, 57, -128, -81, 127, 2, 38, 3, -44, -24, 0, 90, -96, -1, -43, 23, 121, 1, -128, -106, 127, 42, -112, -38, 75, -3, -54, 123, -12, -118, 16, 38, -49, 39, 70, 36, 33, -66, -73, 18, 86, 60, -109, 39, 27, -122, 54, 12, -88, 85, 44, -124, -8, 127, -27, -128, -8, 127, -58, 7, -12, -10, 15, -53, 127, 34, -26, 0, 0, 33, -8, -92, -16, -66, -17, 21, 8, -13, 44, 76, -128, -23, -13, 58, 53, -32, 64, 12, -96, 55, -7, -78, 13, 16, 22, -38, 107, -34, -6, 97, -128, 33, 13, 23, 80, -33, -128, -23, -17, 112, 1, -118, 55, -1, 76, 58, -45, -34, -42, -91, 31, 127, -54, 13, -52, 0, 127, -128, 15, 93, -37, -128, -6, 7, 92, 21, 5, -71, 7, 127, -128, -103, 55, 75, 28, -64, 17, 13, 76, 92, -107, -66, 85, 55, -106, 63, 45, -128, 116, 8, -3, 45, -90, -43, 87, -27, 7, 59, -68, 5, 45, -27, 16, 50, 13, 13, -22, -128, -86, 86, 127, -76, -12, 12, 10, 36, -122, -76, 127, -58, -34, 91, -1, 10, 13, -93, -128, 53, 127, -65, -128, 55, 103, 15, -91, 2, 81, -103, 37, 113, -48, -11, -78, -8, 11, 127, -24, -78, 42, -53, 59, 122, 5, -119, 16, 50, -33, 18, -91, -2, -12, -28, 0, 100, 122, -122, -74, 69, -26, 100, -36, -22, 55, -85, -64, 100, 13, -57, -10, 68, 22, 16, 12, -107, 118, -21, -23, 73, -128, -63, 79, 26, 22, 28, 117, -52, -38, 8, 26, 91, -109, 42, 34, -21, -73, 1, 45, -47, 78, 3, -128, -11, 53, 33, 15, -47, 65, -37, 36, 64, -128, -79, 123, 24, -80, 39, 23, -128, -85, 81, 127, -57, -73, 54, -48, 49, 5, 28, -6, -49, 65, 12, 50, 66, 15, 36, 8, -95, -117, 98, -17, -49, -11, -29, 6, 103, -42, 39, 107, -128, -52, 106, -15, 7, -57, -11, 26, -22, -12, 29, 60, 0, 12, 81, 54, -128, 3, 96, -43, -128, 59, -29, 3, -3, -50, 127, 45, -103, 11, 16, -42, -73, -12, -26, 113, 43, -69, -57, 50, 50, -58, -63, -64, 5, 29, 127, -24, 2, 88, -128, -87, 127, -37, 31, 102, -101, 1, 12, 13, -16, -106, 3, 87, -2, -53, 21, -74, -71, -3, 7, -10, 113, 59, -128, 88, 79, -128, -52, 116, 127, -122, -2, 92, -108, 17, 37, 10, -8, -81, 55, 127, -52, -128, 122, -23, 6, 91, -68, -96, 96, 74, -128, 31, 0, -45, 68, 91, -44, -13, 27, -48, 59, 127, -7, -57, -17, -86, -13, 127, -53, 10, 100, -75, 31, 1, -48, 28, -64, 80, 48, 0, -39, -36, 0, -31, 53, 37, -128, 59, -7, -101, 127, 21, -128, 22, -3, 18, 50, -49, -28, 48, -49, -87, 127, 97, -116, -53, -8, 37, -24, 69, 7, -34, 1, 39, -76, -80, 111, -17, -70, 112, 36, -123, -2, 97, 13, -37, -58, -47, -57, 109, -48, -75, 10, -12, 50, 71, 45, 8, -87, 73, 47, -45, 5, 79, -37, -38, -8, -86, 127, 52, -128, 42, 127, -38, -58, 28, -24, -88, -6, 114, -31, -45, 127, -71, -70, 24, 31, 112, -16, -64, 7, -85, -59, 24, 127, 15, -45, -33, -15, 63, 28, -31, -95, 43, -38, 44, 21, -54, 93, -15, -119, -74, 127, 1, -117, 54, 37, 71, -31, -93, 37, 127, -60, -73, 127, -87, -2, 91, -90, -29, 15, -27, 114, 36, -13, -102, -31, 37, 38, 7, 31, 55, -98, -7, 91, -57, -128, 12, 44, -5, 34, 52, -49, 2, 127, -101, -28, 101, 0, 16, 16, 5, -128, 16, 74, -23, 49, -128, -101, 122, 29, 66, -38, -15, 48, -86, -43, 73, 43, -49, 57, -98, -112, 38, 80, 127, -92, -124, 103, 107, 27, -76, -23, 59, -92, -85, 88, -29, -60, 102, 37, -43, -6, -116, -6, 50, -22, 85, -73, -95, 87, -2, -15, 90, -15, 54, 28, -76, 66, 102, -128, -17, 54, 23, -10, -3, -70, -57, -2, 64, -7, 66, -10, 13, -78, 11, 34, -70, 65, -26, -8, -66, 0, 111, -28, -26, -10, -114, -52, 87, -1, -3, 13, 86, -11, 34, 49, -50, -53, 55, 127, -93, -52, 22, -45, 65, -15, 18, -15, -86, 24, 127, -36, -6, 63, -12, -43, -81, -96, 79, 118, -128, -121, 127, 92, -128, 22, 5, -16, 85, 31, -45, -124, 8, 127, -33, -122, 22, 15, 38, 52, 8, -6, 68, -6, -78, 86, 127, -47, -42, 28, -65, 26, 43, -100, -16, 76, 36, -42, -117, 6, 18, 13, -2, 0, -7, -128, -91, 127, -21, -81, 45, 18, 44, 63, -17, -43, -27, -6, -38, -38, 32, 71, 101, 23, -37, -92, -11, 50, -103, -98, 69, 114, -116, -69, 127, 53, -108, 22, 47, -76, -92, 106, 76, -76, -7, -55, -69, -5, -53, 68, 69, -52, -36, 55, 23, -64, 127, -39, 17, 26, -108, 76, -15, -24, 123, 98, -128, -100, 127, 76, -60, 28, 5, -100, 3, 6, 42, -117, 11, 124, -79, -96, -63, 80, 75, -92, 5, 38, -79, -5, 75, -31, -128, 92, 78, -54, -6, -37, 0, -52, -75, -7, 7, -37, -75, 22, 127, 79, -124, -17, 90, -128, -81, 36, 127, -58, -23, 102, 11, -114, -38, 121, 29, -50, 13, -3, -54, 37, -10, -22, -2, 90, 81, -26, -128, 58, -12, -128, 127, 37, -17, 39, -60, -112, -55, 96, 5, 54, -21, 49, 76, -92, -6, -26, 74, -43, 0, -11, 3, 123, -87, -8, 34, -119, -3, 88, -112, -7, 108, -128, -85, 127, -88, 31, 127, -128, -49, 12, 76, 42, 31, -42, 1, -6, -37, 44, -17, -69, 64, -24, -81, 28, -2, -34, 111, -38, -85, 27, 127, -27, -79, 34, 123, -11, -128, 127, 10, -66, 113, -109, 27, 113, -121, 21, -28, -108, 76, 127, -42, -55, -31, 74, 88, -88, 27, 0, -74, -86, 58, 44, -103, 114, 48, -128, -32, 117, 86, -52, -128, 60, 54, -128, 17, 127, 3, -39, -128, -32, 118, -15, 24, 53, -119, -1, 17, -57, 6, 122, -7, -128, 29, 107, -69, 91, 81, -128, 28, 33, 10, 34, -102, -68, 103, 52, -128, -5, 42, -87, -70, 3, 117, -76, -75, 28, 98, 57, -80, 95, -17, -58, 98, -17, -128, 80, 38, -37, -60, -66, 47, -17, -18, 124, 47, -116, 60, -32, -91, 116, 57, -45, 88, -22, -71, -18, 37, -3, 48, 92, 37, 18, -128, 22, 31, -100, 73, -64, -86, 21, 45, 78, -49, 12, 3, 28, 54, -128, 27, 101, -68, -91, -59, 50, 64, -16, 0, -96, 28, 16, 26, 57, -98, -65, 92, 112, -29, -53, 76, 18, -60, -53, -36, 107, -92, -1, 106, -3, -128, -1, 127, -33, -124, -69, 47, 117, 26, -3, 10, -121, -101, 68, 116, -85, -27, 28, -88, -27, 127, 106, -37, -87, -64, -22, 29, 42, -55, 0, 68, -21, -32, 37, 127, -42, -63, 11, -39, 15, 38, -17, 73, 52, 17, -7, 21, -42, 31, 68, -101, 7, 57, -88, -47, 2, 65, 98, -6, -21, 68, 28, -52, -128, -47, 121, -7, 3, 79, -78, 10, -76, -45, 52, 5, -58, 74, -2, -69, 75, 75, -13, -114, -1, 96, -45, -28, -15, -60, -3, 127, 121, -6, -90, -128, -1, 39, 32, 127, -98, 5, 118, -128, -49, 12, 58, 26, -109, -78, 127, 80, -33, -36, -128, 13, 69, -13, 101, 1, -109, 86, -33, -102, 111, 52, -103, -91, -42, 127, -2, -109, 127, -43, -33, 39, 1, -5, 78, 28, -117, 54, -2, -98, 28, 27, 31, 45, 0, -44, -65, -54, 50, 75, -22, -34, 13, -96, 49, 87, 0, 13, -32, -31, -128, -15, 17, 37, 92, 65, -109, -128, 127, 64, -101, -36, 123, 87, -128, 8, 74, -76, 90, -73, -116, 98, 66, 12, -28, -58, -11, 23, -11, -13, 1, 22, 85, -31, 50, 0, -101, 127, -2, -128, 69, 93, -48, -3, 44, -16, -26, -36, 123, 10, -98, 127, 57, -42, -17, -86, -48, -21, 116, 53, -88, 86, 45, -13, -123, -15, 15, -26, 71, 23, -37, 90, 86, -97, -93, -3, 81, -3, -71, 7, 37, -12, -44, -18, -2, -52, 71, 63, -107, 8, -16, 23, 43, 59, -21, -47, 12, 3, 59, 32, -2, 11, -53, -31, -29, -117, -5, 63, 55, 36, 38, -81, -92, 26, 74, 17, -57, -28, -53, 53, -70, -39, 48, 3, -10, 36, 92, -28, -128, 37, 34, 58, 18, -128, 78, 0, -93, 127, 8, -47, 48, -65, -76, -32, 127, -53, 16, 69, -52, -45, -31, 71, 27, -12, -101, -98, 74, 1, 48, 53, -11, 74, -64, -128, 127, -36, -97, 34, -5, 111, 103, 10, -128, 55, 114, -24, -128, 15, 75, -31, -60, -91, 95, -23, 71, 108, -128, -50, 127, 29, -28, -48, -8, -60, 21, 76, -88, 59, 59, -106, -5, 26, 106, -22, -114, 106, -15, -92, 68, 91, -128, 37, -29, -27, -16, 71, 48, -128, 10, 32, 90, 97, -47, -98, -78, 5, 127, -31, -128, 80, 60, -22, 76, -31, 6, -47, -63, 18, 58, -24, -44, 124, -38, -43, 64, -24, -2, 123, -29, -22, -42, 111, 42, -57, -17, -26, 106, -80, -5, -57, 29, 23, -48, 76, 22, -73, 39, 96, -85, -76, -64, 91, -3, -73, 13, 69, 34, -17, -3, 34, 92, -76, -29, 0, 60, 65, -57, -8, -128, -33, 127, -128, 18, 49, -42, 11, 6, -11, -27, -44, 88, 42, -128, -52, 127, -23, -12, 3, -11, 117, 8, -97, -74, 8, 100, -43, -59, 93, -43, 6, 27, -69, 74, -2, 11, 0, 39, -11, 18, -16, -26, 75, 33, -43, -6, 3, -15, -52, 38, -37, -70, 79, 39, -31, 58, -55, -22, -11, -121, 127, 111, -123, -114, 48, 70, 11, 17, -87, 52, 6, -73, 15, -52, -5, 127, 54, -32, -43, -113, 36, 95, -47, -80, 18, -26, -10, 127, 65, -74, 8, 18, -79, -81, 85, 85, -43, -79, -10, -78, 2, 5, 24, 127, -97, 7, 86, 8, -34, -93, -49, 11, 127, 15, -100, 0, 21, 44, -57, -26, 21, -15, 3, 119, 13, 55, 26, -128, 27, 24, -44, 127, -18, -28, 85, -66, -31, 33, -24, 111, 55, -128, 112, 36, -58, -18, 47, 97, -26, -18, -108, -128, 127, 10, -50, -1, -45, 3, 31, 97, -21, -23, 45, -10, 80, 76, -88, -128, -22, 85, 97, -16, -53, 8, 70, -128, 21, 108, -128, 45, 97, -114, 42, 38, -49, -39, 47, 37, -66, -98, 0, 109, -6, 12, -78, -38, 123, 8, -52, 69, -80, -70, 81, 39, 74, -65, -52, 87, -114, -15, 80, -5, 24, -74, -80, 6, 79, -64, -91, 44, 13, 43, -65, 58, 27, -114, 7, -5, 95, 70, 10, -17, -8, -80, -92, 96, 49, -128, 45, -31, 5, 75, -6, 21, -128, -34, 58, -43, 76, 85, -29, -86, -6, 102, 90, -31, -21, -101, 12, 42, 1, 15, -113, 43, -54, -5, 109, -128, 36, 103, -128, 31, 22, 49, 0, -80, -16, 70, 8, 27, -43, 10, 78, -80, -64, 52, -60, -54, -15, -34, 127, 100, -50, -124, 28, -54, -100, 127, -37, 71, 31, -128, 71, 85, -109, -60, 33, 52, 124, 12, -96, -33, 75, -6, 60, 127, -6, -8, -127, 28, -55, -97, 127, 68, -87, -29, 44, -29, -80, -108, 73, 127, -121, -50, 76, -29, 0, 58, 10, -73, 103, 50, -128, -16, 74, 78, -90, -45, 101, -16, -69, 53, 42, -108, 7, 7, -107, 86, -10, -8, 92, 29, -79, 23, -52, 27, -36, -21, 55, -13, 63, -36, -101, 122, 58, -54, 2, 21, -113, -29, 34, 15, -7, -57, -37, 10, 127, -28, 43, 85, -49, -39, -18, 90, -69, -42, 87, -75, -71, -12, 107, 103, -102, -3, 47, -128, -7, 81, -127, 76, 0, -58, 63, 1, 17, -26, 1, -50, -3, 34, -103, -1, 5, 73, 33, -32, 21, -34, 90, 63, -79, 16, 31, 34, -16, -54, -69, 3, 37, 1, 29, 47, 78, 42, 37, -79, -100, 71, 44, 31, -111, -5, -1, -73, 36, 43, 28, 5, -1, -58, -65, 117, 73, -65, -23, -58, -90, 81, 59, -103, 53, 59, -66, -44, -10, 3, 50, 23, -122, -16, 87, -33, -54, -70, 91, 96, -58, -57, -10, -29, 59, 57, -113, 17, 23, 59, -92, -33, 112, -18, 16, -32, -73, 2, -68, 113, -44, 13, 106, -128, -12, 34, 28, 45, -66, -55, 27, -74, -85, 27, 71, 92, 33, -49, -66, -55, 42, 16, 44, -43, -117, 95, 101, -54, -101, -80, 88, 31, 68, -24, -50, 23, 39, -31, -64, 24, -55, -24, 127, -26, -28, 22, -49, 34, 127, -2, -50, 13, -100, 23, 127, -80, -79, 113, 59, -65, 0, -48, 16, 36, -43, -43, -73, 27, 102, -2, -128, -91, 127, 97, -128, -36, -13, 0, 114, 81, -11, -114, -37, 87, 44, -111, 55, -44, -128, 127, 66, 2, -97, -28, 71, 55, -127, 29, 52, 7, -3, -79, 74, -32, -97, -39, 108, 1, -71, 43, -28, -52, 107, 45, 1, -45, -10, 27, -80, 12, -18, -128, 48, 58, -22, -75, -18, 70, -76, -101, 111, 96, -47, -11, -50, -113, 127, 2, -78, 42, 57, 26, -42, -11, -39, 10, -26, -18, 49, 90, -37, -107, 11, 21, 127, 106, -87, -66, 38, 32, -32, -47, 13, -27, -49, 127, -3, -124, 127, 50, -113, 54, -55, 60, -7, -66, 42, -24, 47, 60, -114, -127, 127, 12, -128, 107, -16, -3, -11, 53, -2, -12, -24, 21, 93, -107, -36, 121, -73, -59, 34, 29, -55, 8, 60, -32, -66, -29, -6, 11, 42, 54, 21, -23, 101, 21, 29, 53, 5, -128, -6, 32, 3, 102, -128, -15, 26, 17, 50, -15, -71, 119, -15, -98, 98, 55, 2, 0, -128, 27, 127, -128, -93, 33, 12, 123, 23, -128, 63, 59, -95, 1, 107, 66, -114, 13, 17, -55, 2, 79, 63, -101, 1, 78, -42, -98, 18, 12, -90, 47, 8, -75, -81, 95, 71, -101, 39, -38, -15, 50, 31, 24, 22, -38, -42, 107, 90, -53, -128, -21, 57, 114, 11, -128, 76, 1, -38, 65, -119, -75, 124, 68, -37, 7, -13, -102, 107, 127, -128, -87, 55, 54, 53, 27, -15, 0, -42, -39, -22, 6, 50, 2, -54, -49, -85, 31, 127, 11, -119, 38, 71, -27, -69, -79, 12, 93, -47, -78, 98, -22, -28, -63, 86, -6, -2, 58, -128, 3, 27, 33, -17, -54, 69, 103, 8, -44, -42, 23, 0, 34, 10, 102, -22, -27, -8, 22, 33, -24, -66, -1, -15, 79, 48, 15, 63, -128, -37, -45, 48, 106, -64, 0, 17, -5, -74, -87, -17, 59, 50, -50, -102, 116, 18, -93, 55, 42, -80, -44, 48, 28, 66, -18, 76, 106, -128, 26, 2, -21, -49, -81, 116, 60, 52, -64, -57, 8, 26, 57, -128, -34, 37, -31, 26, 69, 11, 52, -87, -16, -22, -26, 127, -8, -57, 48, -38, -17, 23, -5, -69, 3, -98, -91, 97, 127, -17, -128, 26, 38, 75, 12, -26, -81, 33, -29, 16, 34, -114, -15, 28, 38, 71, 124, 18, -128, 57, 11, 16, 50, -128, 0, 64, -49, 23, 127, -95, -109, 2, 109, 45, 48, -53, -96, 15, -7, 50, 127, -24, -93, 102, -26, -64, -2, -16, -11, 31, -10, 29, 17, 50, 37, -12, -81, 38, 0, -87, -22, 68, 29, 32, 103, -119, 29, -22, -91, 127, -2, -119, -2, 122, -68, 1, 24, -39, -47, 44, -37, -26, 44, 10, -6, 114, -31, -57, 122, -21, -8, 45, 13, 10, -97, 3, -54, -54, 127, -10, -96, 18, 66, 36, -75, 49, 6, -17, -21, -7, -5, -27, -66, 49, 119, -107, -33, 118, -7, -111, -16, 12, 114, 113, -6, -128, -16, 127, -79, -55, -11, 22, 76, 23, -117, -113, 106, 66, 2, -114, -55, 28, 33, 11, -118, 17, 103, -16, -60, -38, 69, 33, -57, 6, 31, -33, 44, -16, -54, 127, 38, -100, 8, 2, -44, 69, 24, -128, 22, 59, -52, -65, -45, 12, 123, -48, 0, 28, -13, -92, 18, 23, -26, -68, 60, -26, -70, 75, -32, 29, 18, 58, -78, -107, 93, 74, -66, -36, 127, 91, -128, -32, 55, -43, 114, -38, -38, 85, 18, -65, -128, 95, -29, 5, 127, -18, -29, -108, -58, -32, 100, 97, -128, -93, 22, 100, 96, -97, 50, 52, -128, 96, -31, -53, 42, -73, 103, 117, -21, -50, -86, 52, -8, -85, 48, -5, -52, 27, 64, 2, -34, -11, -34, -7, 7, -44, -88, -10, -90, -3, 52, -32, 37, 28, 47, 27, -53, -24, 28, -23, -66, 127, -23, -45, 27, 54, -85, 6, 52, 11, 0, -118, 49, -5, -96, 91, -38, 13, 26, -98, -18, 90, 3, -12, -57, -63, 45, 64, 26, 23, 7, -49, -8, -128, -44, 48, -63, 69, 3, 21, 49, 33, -107, -34, 59, -3, 1, 50, -18, 38, 91, -71, -49, -18, -53, 69, 31, -38, -42, -55, 34, -1, -75, 34, 45, 12, -128, 34, 50, -98, 24, 127, -95, -49, 65, -23, 80, 15, 16, -117, -58, 127, 8, -128, -16, 6, -38, 24, 127, 31, -63, 3, -85, -87, 50, 127, 39, -114, -2, -42, 6, -7, -65, 112, 55, -29, -90, 22, 36, -60, 85, 113, -119, -39, 127, -22, -64, -66, 53, 49, -2, -17, -79, -55, 70, 86, 50, -64, -128, 79, 70, -18, 17, -5, -87, -38, -5, 0, 98, -21, -70, 5, -44, 27, -66, -8, 36, 44, 36, 58, -80, -79, 71, 13, 0, -53, -13, 80, 57, -22, -34, -5, 127, 97, -42, -111, -55, -15, 90, -10, -5, 6, -128, 1, 44, -29, 108, 28, 3, -32, -45, 122, 1, -5, -60, 32, 74, -109, -60, -1, 65, 15, -37, 42, -1, -49, 111, 55, -98, 21, -66, -50, 37, -29, 64, 29, -70, -26, 113, -97, -27, 33, 53, -34, -108, 44, 6, 127, 49, -87, -33, -18, 127, 42, -7, -70, 44, 69, 15, -63, -43, -18, 60, 109, -80, -50, 3, 44, 57, -102, 0, 0, -34, 22, -26, -7, 13, -28, -38, -70, 81, 39, -123, 31, -52, 66, 74, -38, -38, -43, 96, 29, -95, -18, 23, -124, -38, 37, 118, -33, -29, 86, -3, -76, -26, 21, -53, -1, 127, 18, -103, 74, -74, -7, 54, -96, 48, -24, 60, 123, -101, -17, 36, -128, -7, 71, -91, 66, 79, -128, -81, 79, 113, 27, -28, -91, -86, 114, 42, -114, 0, 127, 74, -108, -48, -5, 15, -52, 0, 68, -65, -49, 79, -16, 3, 18, 65, 69, -112, 8, 117, -76, 57, 31, 1, -1, -27, -95, -22, 44, -31, 112, -15, -71, 34, 112, 36, 0, 48, -128, -45, 12, -12, 127, -54, -39, 127, 0, -128, -88, 39, 127, -29, -98, 63, 1, 75, 127, -123, -123, 58, 42, 102, -8, -59, 108, 70, -32, -70, 5, -122, -87, 29, 59, 8, -12, 127, -70, 36, -1, -128, 45, 127, -22, -81, 17, 10, 127, -50, -80, 127, -44, -48, 66, -22, 47, -23, -65, 65, -63, -49, 121, -34, -50, -13, 3, 91, -57, -11, 97, -49, -5, 92, 71, -58, -1, -108, 2, 117, -128, -88, 122, 24, 0, -28, 54, 13, -22, -21, -74, 112, 64, -128, -37, 43, 8, 80, 81, -78, 57, -17, -76, 18, 106, -34, -6, 70, -112, -12, 31, -39, 32, -64, 36, 1, -60, 59, 47, -117, 49, 109, -36, -63, -128, -44, 127, -33, 3, 43, -59, 29, 34, -1, 18, -36, -128, 65, 44, -65, 21, -79, 112, 1, -113, 117, 12, -17, -18, -73, 81, 0, -100, 98, -53, -59, 2, 116, 39, -22, -38, 32, -1, -128, 80, 28, 0, 64, -102, -68, 27, 95, -11, -78, 127, 31, -128, 27, 44, -2, 91, -92, 47, -21, -128, 24, 96, -8, 88, 107, -44, -128, 23, -13, -70, 53, 44, -79, -36, 127, -33, -38, 37, -13, 36, -31, -119, 96, -54, -43, 60, 43, 21, -88, -113, 92, 50, -68, 71, -37, -75, 58, 29, -81, -92, -7, 127, 68, -119, -66, 73, 43, 28, -87, -86, 97, 58, -68, -24, 54, -123, -98, 127, -91, 10, -11, 33, 31, -49, 73, 24, -128, -1, 87, -42, 21, 47, -71, -24, -39, 58, -2, 33, 57, -58, -60, 18, 31, 66, -34, -69, 127, 1, -128, 106, -16, -118, 107, 22, -10, -15, -87, 70, -69, 29, -2, -16, 47, -43, -73, 36, -13, -45, 38, 52, 29, -52, -103, -52, 45, 36, 11, -7, -97, 95, 43, -85, -32, 13, -7, -33, 127, 17, 3, -70, -64, 31, 109, -68, 17, 2, 0, -26, -10, 28, -109, 70, -10, -13, -33, 65, -8, 8, 24, -74, 73, 78, -22, 7, -103, 0, 127, -127, -96, 127, -18, -23, 0, -47, 127, -32, -11, 95, -27, -33, -31, 80, -15, -11, 34, -17, 22, 36, 127, -2, -47, 21, -37, -16, 39, 33, 96, 119, -123, -8, 87, -92, -65, 97, -2, 7, 53, -128, -11, 55, -49, 69, 86, -97, 26, 91, -128, -128, 11, 28, 45, 78, 0, -23, 28, 8, 0, -50, -5, 96, -92, -54, 34, 39, -10, 64, 37, -114, 91, -26, -24, 7, 74, 28, -57, 92, -36, 12, 78, -75, 32, -73, 54, 1, -65, 53, 42, -97, 33, 3, 7, 76, -80, -128, -16, 107, 44, -29, -16, -60, -5, -74, -21, 37, -33, 76, -88, -18, 59, 22, -107, -42, 1, -38, 127, 50, -16, -18, 5, -13, 15, 3, -71, -32, 69, -121, -63, 127, 45, -112, -50, 71, 11, -106, -24, 28, -16, 64, 124, 11, -91, -96, 0, 90, -21, 106, -57, 12, 53, -18, -10, -65, 34, -52, -66, 117, 3, 3, 42, 80, 27, -38, -22, -73, -113, 127, 69, -128, 15, 58, 48, 39, -66, -128, -5, 109, 92, -95, -54, 29, -63, -54, 127, 88, -128, 64, 3, -106, 37, 79, -31, -69, 70, 121, -28, -71, 71, -95, -12, 36, -2, 23, -57, -37, 73, 50, 37, -31, 7, -26, -128, -22, 95, 122, 11, -75, 7, -117, 37, -5, -5, -24, -43, 33, 107, 63, -69, -17, 21, -95, -118, 48, 108, -59, -21, 3, -123, 69, -16, 81, -7, -122, 27, 118, -31, 73, 8, 6, -53, -87, 33, 117, 1, -39, -26, -6, 54, 102, -57, -58, 38, 1, 127, -70, -5, 73, -55, 26, -75, -21, 78, -73, -7, 75, -128, 10, 118, -113, -11, 71, -64, -8, -7, -10, -80, -2, -48, 5, 68, -74, -86, 118, 81, -128, -66, 108, 92, 10, -64, -98, 42, 23, 24, 1, -55, 90, -16, -73, 6, 127, -52, -24, 127, -29, -45, -90, -1, 102, -116, -69, 58, -1, -3, 127, -24, -103, 81, -47, -59, 127, -31, -48, 21, 23, 90, -65, -63, -64, 57, 79, -116, 57, 22, 42, 16, -128, 5, 24, 122, 5, -75, -16, 33, 75, -86, 39, 109, -53, -16, -128, 5, 127, -63, -2, -3, -90, -16, -55, 44, -11, 32, 64, 13, -121, -7, 63, -101, 113, 55, -128, -16, 127, -58, -12, 55, -92, 15, 29, -93, 7, 78, 45, -39, -97, 96, -34, 10, 26, -59, 23, 24, 109, 57, -128, -127, 81, 102, -92, -2, 23, -49, 116, -15, -57, 69, 50, 6, -113, -53, 111, 10, -5, -17, -128, -50, 87, -1, 74, 59, -73, -76, -28, 88, -7, 10, 75, 42, -86, 36, 7, -50, 122, 70, -76, -113, 24, 24, -96, 91, 108, -128, -11, 127, -24, -22, -117, -73, 127, 73, -43, -97, 27, 60, -39, -128, -42, 65, 60, 7, -116, 101, 93, -23, -5, -100, -86, 31, 103, -44, -75, 74, -7, -121, 71, -2, 34, 70, -108, 31, 28, -100, -33, 90, -26, 101, 45, -100, -8, -26, 107, 8, -124, 81, 15, 69, -68, -36, 69, 44, 52, -36, -55, -92, 60, -34, -63, 86, -121, 48, 65, -58, -80, 39, 127, -128, -33, 75, -42, 70, 16, -113, -54, 92, 86, -69, -36, 69, -118, -102, 127, 113, -3, -109, -95, 90, 31, -21, -44, -37, 16, -114, -65, 113, 60, -121, 26, -2, -12, -24, -68, 34, 37, 11, -69, 8, -24, 92, 24, -128, 127, -26, -128, 127, 39, -95, 63, -42, -63, 49, -48, -33, 113, 18, -119, 38, 119, -124, -100, 127, 26, -31, -23, -48, 11, 81, 73, -44, -22, 127, -21, -96, 127, 0, -122, 39, 124, -112, 28, 29, -29, -50, 26, 50, -18, 60, -108, -36, 127, -70, -97, 27, 96, -7, -73, 76, 43, -29, 21, -128, -12, 31, -54, 69, 39, -21, -88, 29, 86, -112, 92, 23, -128, 87, 87, 3, -69, 31, -42, -68, -6, 36, 95, -111, -86, 50, 127, 93, -128, 31, 127, -54, -128, -34, 44, 81, 55, -74, -63, 6, 32, -23, 42, 36, 29, -48, -71, 13, -5, 60, 58, -44, -76, 17, 42, -47, 38, 8, -90, 81, 8, -91, 57, 50, -11, 71, -42, -70, 27, 70, 49, 7, 34, -85, -68, 98, 43, -26, 59, 27, -128, 5, 12, -18, -27, 65, 68, -17, -101, -128, 96, 87, -92, -65, 127, 28, -24, -71, -8, 127, -32, -128, 32, 33, -43, 78, 79, -7, -124, 24, 48, -66, -18, 93, -118, -15, 127, -18, -44, -128, 60, -1, -32, 106, -98, -39, 18, -92, 86, -21, -90, 85, 17, 58, 64, -33, -38, 29, -11, 33, 3, 68, -64, 15, 127, -128, -8, 102, 45, -107, 3, 76, -75, -37, 24, 44, -112, -91, -15, 127, 2, -128, 34, 52, 57, 49, -11, 7, -117, 27, 10, -79, 64, -22, -73, 37, 22, 52, -55, -45, -1, -21, 42, 98, 74, -128, 7, 127, -108, -37, 114, -73, -17, -66, 31, 28, -128, 71, 48, -73, 48, 69, 1, -85, -68, -39, 127, 69, -18, -103, -112, 127, -8, -101, 75, 96, -74, -113, 122, 36, -128, 102, -5, -2, 2, -109, 57, 26, 78, 53, -57, -49, 8, -24, 42, 55, -97, -2, 10, -86, 70, 33, -109, -74, 127, 103, -128, -55, 43, -43, 127, -3, -128, 37, 23, 38, 43, 28, 54, -53, -31, 27, 73, 92, -26, -59, 11, 96, -95, -113, 59, -12, 100, 66, -121, 54, 34, -78, -53, 91, 32, -117, 118, 28, -109, -57, 102, 69, -58, -38, 47, 43, -43, -54, 0, 127, 0, -17, 23, -43, -128, -70, 127, 73, -33, -128, 12, 32, -58, 95, -96, 27, -31, -114, 90, 36, -34, -27, 127, 38, -101, 7, -50, 54, 68, -81, 5, -47, -47, 60, -80, 8, -38, -76, 127, -64, -34, 96, 0, -106, 33, 124, -128, 33, -21, -8, 37, -47, 119, -39, 43, -11, -1, -17, -93, 97, 98, -118, -86, 102, -45, 29, 58, -75, 111, -24, -88, 43, 80, 48, -93, -60, 36, -2, -79, 45, -43, -8, -31, 87, 85, -18, -103, -31, -5, 2, 33, -64, 81, 63, -12, 26, -81, -91, 127, -23, -85, 50, 49, -12, -34, -10, 122, -49, 16, 10, 5, 109, -49, -36, 17, -79, -3, -73, 64, 103, -102, -98, 92, -49, -2, 44, 6, -117, -12, 127, -111, -109, 38, 127, -7, -47, 117, -86, -45, 102, -42, -49, 54, 106, 47, -124, -90, 74, 0, -55, 22, 97, -17, -85, -68, 28, -6, -49, 91, 95, 42, -50, -24, -93, -26, -2, 55, 36, -76, 127, 88, -128, -81, 27, 27, -22, 80, 52, 18, -95, -118, 96, 11, 38, 127, -87, -107, -15, 59, 98, 45, -73, -66, 50, 8, 17, 16, -128, 88, 98, -128, 59, 0, -66, 36, 36, 43, 87, -87, -70, 127, -91, -6, 3, 2, 88, -70, 31, 17, -21, -47, -48, -64, 81, -48, -22, 70, -18, 2, -38, -57, 36, -29, -26, -60, 15, 127, -47, -95, 92, 36, -123, 53, 0, -88, 47, -48, -107, 111, -17, 69, 10, -34, -3, -60, 114, 88, -22, -85, -23, -7, -111, 22, 127, -21, -68, -22, 10, -86, 79, 50, -16, -53, -28, 11, 55, -33, -24, 86, 22, -53, -21, -80, -58, 127, -7, -128, 124, 0, -28, 47, 2, 15, -128, 24, 26, 2, -49, 45, 73, -128, -15, 88, -44, 66, 69, -128, -80, 75, 118, -91, -114, 127, 3, -36, 59, 27, -24, -33, 79, -65, -123, 114, 127, -113, -57, 38, -79, 90, 33, 3, 55, -12, -86, -101, 107, -3, -68, -27, 101, 17, -108, 122, 95, -113, -92, 38, -53, 79, -24, -109, 45, 27, 127, -43, -32, 49, 5, 22, 90, 28, -128, 31, 47, -36, -101, -1, 127, -54, -60, 57, -3, -12, -16, -23, -74, -76, 26, 68, -49, 10, 96, -54, 27, 36, -68, 127, 36, -73, -23, 10, -11, 23, 10, -101, 16, 88, 31, -47, 86, -38, -124, 113, 123, -5, -109, -65, -53, 95, 118, -128, -73, 76, 7, 69, 63, -69, 22, -34, 53, 113, -55, -128, 21, -12, -58, 127, 22, -36, -71, -27, 121, -59, -114, 127, -33, -24, 10, -55, 36, 127, -54, -68, 18, 3, -28, 93, 69, -37, -121, 8, 107, 0, 10, -91, 38, -58, -73, 92, 80, -29, 32, 3, -37, -92, -21, 124, -2, -39, -111, -80, 127, 11, -12, -69, 47, 93, -6, -58, -79, 92, -79, -111, 124, 108, -65, -54, 79, -2, 5, -13, -128, 91, 0, 8, -52, 7, 103, -24, -43, -128, -53, 97, 45, 47, -2, -81, 24, 18, 34, 79, -107, -12, 108, -12, -81, -73, -16, 6, 121, -63, 22, -37, -109, 52, 127, -26, -128, 127, -18, -2, 112, -107, -85, 22, 127, 27, -91, -32, 100, -65, -87, 23, 119, -32, 42, 3, -74, -5, 43, 15, -37, 33, -11, -10, 55, -58, -5, 75, -128, 26, 63, -128, -48, 127, -3, -108, 47, 102, -3, -70, 68, 43, -76, -10, 63, -44, -128, 18, 127, 15, 3, -90, -63, 23, 98, -57, -3, 79, -117, -92, 117, 123, -128, 36, 80, -114, 87, -68, -128, 114, 37, 76, -60, 11, 55, -128, -1, 92, 21, -73, -6, 55, 13, 44, 48, -86, 38, 12, 5, 57, -111, -53, 45, -31, -47, -27, 71, -12, -86, 80, 47, -57, -16, -128, 6, 48, -86, 121, 90, -74, -128, -52, 127, 0, -37, 31, -33, -8, -92, 23, 58, -2, -59, -28, -3, 68, 76, -128, -59, 44, -16, 17, -2, 127, 5, -26, -6, -27, 85, -53, -70, 127, 27, -91, 15, 21, 118, 97, -39, 15, -54, -97, 43, 59, -10, 7, -48, -47, -91, 68, 112, -128, -111, 127, -29, -73, 102, -27, 54, -31, -49, 119, 45, -52, -1, 31, -42, -59, 12, -29, -11, -29, 70, -18, 59, 27, 17, -17, 10, -81, -86, 127, -45, -58, 96, -44, 22, -18, -18, 47, -42, 87, -52, 54, 2, -23, 55, -7, -95, -65, -6, 70, 16, 10, 37, -98, -74, 90, 80, -117, 36, -34, 48, 127, -128, -32, -31, -71, 123, 63, -55, -97, 12, 111, -93, 48, 54, -5, 8, -7, -102, 32, 29, -52, 32, -87, 47, 71, -27, -49, -128, 39, 113, -128, 32, 15, 2, 116, -87, -49, 42, 54, -31, 26, -32, -71, 43, 52, -90, -80, 74, 6, -78, -28, 5, -33, 81, 0, 69, 21, -16, -98, -71, 127, -60, 74, 91, -69, 11, -112, -66, 65, 121, 36, -106, -26, 13, -29, 34, 103, 22, -87, -24, 127, -1, -50, -69, -54, 127, 114, -64, -68, 47, 18, -128, -128, 127, 127, -60, -78, 47, 5, -43, -7, -71, -97, -23, 121, -12, -18, 24, 42, 27, -29, 6, -88, -50, 114, -6, -102, 92, 127, -33, -57, 11, 22, -52, -58, 36, -63, -108, 116, -24, -121, 118, 78, -103, 60, 0, -63, 8, 57, -31, -98, 55, 127, -71, -24, 66, -47, 28, -37, -34, 26, 102, -54, -86, 80, 81, -101, 48, -33, -122, 53, 22, 112, 80, -91, -3, -52, 43, 119, -26, -128, -95, 60, 127, -50, 3, 32, -47, 2, 5, 52, 0, -69, -117, -33, 42, -22, 60, 37, -47, 75, 39, -33, 8, -12, 71, 119, -98, -59, 123, -93, -48, 127, -63, -60, -22, -24, 127, 44, -53, -23, -15, -1, -81, 43, 76, -93, 8, -57, -23, 98, -11, -128, -50, 27, 3, 127, -70, -39, 64, 60, 0, -15, 7, -8, -109, 16, -45, -97, 95, 76, 13, -121, -37, -13, -44, 49, 90, -88, 22, 55, -127, 39, 73, -63, 16, 66, -103, -1, -5, -7, 48, -128, 27, 90, -119, -49, 118, 11, -10, 12, -24, 34, 70, 50, -31, 13, -76, -55, -18, -22, 10, 29, 127, 31, -42, -26, -13, -95, 1, -10, 95, 0, -121, 91, 100, -102, 8, 17, -37, -32, 43, 73, -27, -63, 7, -7, -34, 109, 49, -88, -112, 92, 100, -128, 6, 90, -5, -59, 24, -33, -38, 90, -23, -2, -16, -58, 113, -58, -7, 42, -59, 23, -38, 108, 75, -60, -76, -74, 98, -16, 12, 102, 42, -85, -22, 38, -128, 2, 127, 7, -60, -58, -15, -32, -52, 127, 22, 7, 73, -128, -63, 42, 37, 31, -47, 0, 0, 50, 39, 47, 2, 44, -27, -69, 11, -39, 127, -3, -68, 108, 55, -128, -88, 70, 1, -3, -3, 75, -6, -87, 112, 43, -75, -48, 107, 11, -78, -92, 96, 97, -74, -76, 6, 95, -32, -32, 43, -63, -128, 26, 74, -85, 60, 102, -44, -113, -38, 127, 78, -100, 50, 11, -128, 6, 127, 50, -10, -116, -128, 127, -6, -31, 5, 31, 31, 2, -11, -59, -26, 34, -87, 57, 86, -54, -15, -95, 28, 79, -128, -6, 33, -59, 15, 39, 81, -38, -21, 102, 22, -39, 18, 45, 64, -5, -100, -16, 49, -79, -45, 32, 127, -17, 59, 18, -22, 12, -43, -2, -60, 31, -59, -16, 108, -97, 11, -7, -87, -38, 106, 71, -112, -52, 2, 5, -47, 80, 101, -48, -28, 22, -24, -73, -111, 66, 124, 2, -117, -33, 31, 17, -32, -128, 50, 86, -64, 32, -78, 47, 127, -128, 3, 47, -24, -43, 63, 63, 5, -11, -101, 28, 42, -95, -32, 109, 108, -108, -2, 21, 55, -2, -96, 54, 6, 92, -76, -3, 93, -127, 32, 65, -76, -13, 124, 31, -91, 10, -17, -31, 7, 55, 113, -1, -69, 69, -70, -98, 127, 39, -108, 37, -98, 13, 39, -58, 75, -5, -73, 11, 66, 73, 26, -42, 48, -26, -124, -8, 127, -28, -70, -27, 78, 8, 0, 0, -76, 127, 36, -116, 32, 127, 36, -96, -33, -55, 64, -8, -52, 127, -48, 2, 1, 28, -48, -85, 32, 2, 39, -23, 26, -59, -18, 74, -18, -50, 85, 37, 24, 91, -88, -119, 103, -17, -15, 15, -44, 16, 16, 57, -74, 18, 28, -42, 37, -128, -74, 81, 26, 80, 27, -128, 71, -24, -38, 21, -44, 12, 70, 127, -116, 34, -11, 17, -13, 1, 3, -28, -10, 52, -2, -54, 63, -109, -44, 112, -86, 13, -23, -6, 66, 13, 2, -79, 42, -66, -27, -32, -22, 32, -52, 79, 13, -32, 68, 31, -60, 103, -28, -42, 127, -1, -109, 31, 88, -16, -53, -113, 28, 100, 13, -102, -1, 49, 15, -11, 12, -42, -13, -39, 0, 68, -11, 5, -128, -57, 68, -6, -6, 49, 86, 66, 16, -32, -76, -7, 0, -122, 76, -22, 7, 59, -93, -2, -24, -24, 15, 0, 109, 117, -71, -66, 69, -31, -50, 103, 23, -33, 64, -12, 5, -26, -60, 75, -49, 57, 13, -16, -74, -43, -7, 112, 127, -128, -69, -28, 38, 59, -59, -27, 42, 64, 17, 58, 1, -43, -33, 76, -87, -107, 95, 96, -16, 1, -26, -15, 28, 17, -65, -12, -54, -43, 88, -79, 42, -33, -78, 49, 37, -3, -29, 69, -117, -128, 127, 60, -33, -70, 3, 75, -39, -98, 34, 127, 17, -22, -53, -66, 48, -90, -49, 2, 65, -13, -45, 76, -16, -128, -7, 52, 58, -70, -32, 127, -60, -69, 68, 101, -26, 42, -21, -15, -88, 44, 92, -36, 11, -98, -52, 70, 10, -128, -58, 108, 28, 28, -12, -123, 93, 92, -102, -44, 52, 21, -123, 43, -80, -23, 113, -75, 6, -43, -59, 118, -50, 63, 48, -6, -45, -128, 118, -24, -74, 5, 93, 91, 2, -118, 17, 87, -128, -29, 71, -75, 0, 127, -86, -49, 92, 37, 29, -119, 45, -59, 29, -13, -128, 127, -10, -2, 109, 53, -38, -128, 112, 22, -42, 85, -64, -33, 13, -5, -97, -69, 116, 37, -128, 81, -42, -16, 90, 18, -128, 0, -8, 59, 100, -128, -3, 121, -22, -95, 58, -29, -59, 118, 23, -114, 65, -7, 48, 27, 15, -78, -10, 101, -29, 3, -33, -21, -23, -80, 28, 27, -128, 49, 57, -22, 29, -128, -16, 38, -39, -10, 18, 53, -92, -92, 127, 90, -128, 10, 1, -85, 109, 107, -12, -98, -3, 2, -90, 2, -45, -27, 39, 17, -7, -36, 48, 31, 15, -18, 81, 111, -63, -74, 28, 43, -29, -29, -2, 55, -71, 8, 109, 5, -60, -18, -39, -34, -5, 68, -86, -18, 7, -11, -31, 8, 87, -34, 8, 70, -65, -86, 65, -98, 37, 43, -22, -23, 44, -34, -124, 127, 87, -47, 0, -91, -13, -10, -96, 10, 68, -2, 106, 23, -26, -103, -80, 91, 36, 64, -36, -128, 29, 38, -39, 15, 93, 70, -37, -59, 65, -5, -88, 36, 0, -55, -21, -3, 109, -1, -24, -21, 45, 48, 33, -11, -44, 88, 45, -128, 36, 39, -128, 15, 92, -33, 1, 7, -76, -5, 124, 102, -42, -128, 24, -10, -18, 118, -47, -88, -18, 127, 3, -5, -23, 91, -49, -36, 127, 6, -64, -11, -87, 26, -27, -128, 23, 127, -8, -87, -31, 0, 47, 103, -23, 17, 59, -54, -38, -101, -112, 127, -27, -75, 100, -17, -15, 59, 100, -66, -47, 88, -69, 63, 63, -87, 66, 54, -113, -55, 0, 32, 57, 15, -60, 86, 24, -128, 81, -2, -59, 107, -86, -33, 0, 23, 80, -48, -92, 45, 81, -23, 81, 2, -128, 10, 127, -102, -68, 53, 16, 45, 33, 65, -128, 24, 119, -76, -122, 47, 118, -45, -44, -81, -49, 127, 55, 0, -117, 15, 13, -1, -16, -37, 32, 18, 109, -50, -50, 127, -49, -43, 23, 34, -8, -78, 50, -24, -127, 127, -29, 22, 48, -44, -91, 29, 54, -1, -1, -28, -16, 43, -60, -23, 127, -81, -12, 50, -80, -74, 69, 66, 15, -103, -10, 37, 13, -11, 23, 45, -106, 44, 37, -23, -28, -21, -2, -111, 27, 3, 37, 127, -2, -33, -75, 23, -64, -58, 86, 31, 1, -43, -16, 49, 29, 87, 34, 12, 63, -117, -53, 8, -39, 15, -2, 108, 109, -58, -12, -59, -1, 13, -70, 47, -8, 50, 17, -64, 127, 50, -42, -66, 38, 75, -69, 59, -34, 17, 64, -108, -45, 18, 78, 27, -15, 44, 124, -86, -128, 127, 29, -15, 107, -70, 0, 64, -28, -128, -114, 127, 69, -42, 31, -66, -79, -6, 127, -1, -17, 34, -78, 69, 3, -8, -100, 38, 2, 34, 91, -128, 0, -12, 45, 53, -53, 32, -15, -49, 50, 3, -119, 5, -5, 91, 53, -128, 71, 26, -88, 43, -95, 50, 60, -57, 8, -7, -48, 44, 16, -116, 107, -32, -98, 121, 29, 3, -42, -101, 5, 17, 81, 1, -5, -101, -22, 79, -42, 17, -50, 90, 10, -114, 109, 80, -13, -79, -39, -12, -23, 127, 5, -116, -13, 107, 119, -13, -65, -58, 81, 54, -70, -11, -57, -45, 86, -112, -102, 74, 86, -17, -55, 127, 2, 18, 10, 38, -91, 1, -3, -85, 124, 11, -63, 57, 109, -122, -70, 74, 16, -17, -5, -1, -18, 114, 87, -128, 32, 121, -112, -78, 127, -32, 16, -39, -128, 80, 8, -17, 31, 13, 31, 106, -2, -42, -12, -29, 33, 49, -128, -60, 63, 15, 49, 10, -47, 1, 53, 122, -97, -5, 32, -100, 11, 60, 36, 0, 91, 13, -49, 91, 0, -27, 17, -119, -16, 13, 47, -12, -91, 91, 38, -58, -69, -45, 127, -1, -75, 26, -15, 45, -31, 27, 80, -70, 58, 87, -80, -26, -32, 88, 11, -2, 48, -106, -69, 42, 90, 92, -22, -11, 5, -98, -39, 114, -7, -90, -23, 114, 50, -70, -37, 50, 93, -8, -29, -24, -55, 87, 60, -122, -2, -38, -71, 55, 31, -27, 47, 111, -113, -91, 127, 69, -74, 55, -13, -31, -63, -6, 49, 0, 55, -18, -127, 33, 1, 39, -42, -23, 118, -117, -93, 127, 18, -52, 127, 21, -91, 0, -2, -6, 44, -71, -50, 22, -3, 111, 107, -98, -73, 21, 121, -68, 32, -36, -2, 2, 34, -75, 10, 123, -128, 73, 29, -111, 10, 2, 111, 32, -27, -68, -88, 48, 34, -24, 17, 18, -91, -8, 121, -49, -18, 43, -66, 1, -128, -15, 36, -81, 103, -2, 49, 78, -128, -53, 127, -1, -81, 101, -81, -57, 42, 5, 106, 24, -28, -53, -66, -68, -31, 63, 79, -85, -28, 65, -71, 38, -3, -23, 92, 47, -37, -33, -7, 31, 47, -59, 80, -45, -96, 28, 71, 60, 5, 0, -26, 27, -43, 85, 74, -108, -28, 17, 27, -91, -73, 127, 64, -109, -47, 21, 127, 28, -43, -69, 114, -28, -98, 127, -64, -57, 127, -23, -5, -29, -128, -1, 127, -45, -117, 114, 44, -10, -64, -63, 97, -1, -108, 24, 88, -38, 13, 26, 21, 107, -73, -42, -57, 45, 70, -92, -22, 55, 103, -79, 36, 100, -113, 13, 86, -73, -68, 15, -52, 43, 88, -128, -93, 127, -11, -36, -58, 53, -39, -5, 127, -85, -78, 102, -68, 1, 127, -122, -118, 114, 15, -112, 57, 101, 38, -52, -87, 22, -27, 58, 13, 70, 39, -111, 71, -87, -96, 23, 127, -22, -11, 75, -53, -102, 22, 74, 34, -49, 3, -93, -70, 52, -26, 101, 102, 1, -128, -98, 54, 18, 74, 37, -87, 1, -17, -2, 93, 0, -8, 38, 28, -32, -18, 5, 39, 117, 48, -101, -48, 86, -15, -5, 87, -52, -80, 73, -18, -32, 90, -15, -22, -11, -93, -78, 127, 2, -113, 60, 32, 11, 49, 31, -52, -1, 26, -128, 0, 108, -91, -79, 36, 92, 49, -74, -75, 0, 127, 17, -65, 66, 53, -98, -79, -6, 21, 33, 5, 43, 44, 28, -122, -18, 92, 23, -52, -36, 54, -81, -64, -3, 12, 87, 54, -128, 43, 116, -128, 42, 0, -11, 78, -103, 87, 113, -128, -69, 11, 60, 90, 26, -87, -128, 58, 15, 74, -44, 8, 98, -97, -86, 103, 52, -29, -37, -28, 1, -79, 23, -7, -48, 0, -86, 64, 33, 37, 58, -65, -128, 5, 74, -90, 96, 43, -59, -64, -16, 113, -87, -53, 47, 24, -1, 127, -34, -8, 70, -1, -100, -39, 21, 48, -93, -32, 85, -26, -5, 5, -59, 44, 127, -36, -53, 44, -108, -63, -8, 73, -1, -86, 127, -5, -69, -24, -8, 114, -66, -73, 127, 10, 18, -32, -73, 127, 48, -22, -76, -70, 13, 37, 109, -55, -112, 108, -1, -21, -7, 18, 18, 0, 91, -43, 45, -8, -57, 127, 50, -128, -79, 58, 74, 54, -26, -10, 2, -92, -1, 102, -48, -16, -33, -53, -42, 50, 0, -33, 127, -59, -23, -11, -7, 34, -23, 5, 34, 73, -42, 119, 74, -128, 1, 12, 100, 91, -27, -74, -117, 22, 37, 32, -45, 34, -52, -57, 54, -42, 64, 1, -49, 7, 0, 75, -7, -54, 50, -3, -11, -1, -60, -73, 64, -114, -28, 127, 7, -66, -76, -54, -11, -7, -11, 118, 127, -97, -118, 60, 58, 59, 10, 0, -108, -103, 108, 59, -22, -38, -57, 15, -8, -90, -26, 64, -3, -86, 60, 33, 44, -68, -8, 127, -128, -33, 87, 44, 5, -60, -69, -49, 50, -27, -39, 122, 3, -128, 66, 11, 26, -22, -107, 47, 65, 2, -86, -73, 116, 91, -70, -36, 53, 74, -90, -22, 10, 28, 11, -119, 18, -45, 27, 17, -43, -22, -15, 127, -18, -128, 55, 36, 7, 65, 53, -102, -65, 127, -60, 17, 58, -79, -28, -22, 26, 78, -97, 68, 76, -52, -60, -58, 119, -87, -7, 43, -78, -33, 45, 100, -66, 50, 107, -68, -59, 24, 26, 7, -26, 15, 15, -103, -31, 127, -11, -34, 45, -55, 21, -11, -78, 127, 64, -128, -64, 87, 63, -27, 0, 78, 39, -76, -47, 11, 52, 27, -128, -34, 66, 8, -48, -70, 106, 32, 39, 60, -12, -91, -111, 38, 73, -52, -22, 2, -11, 27, 58, -128, -114, 91, 127, 42, -17, -96, -59, 86, -57, -21, -1, 39, -42, -39, 107, 8, -16, -29, -42, 21, -91, -121, 92, -5, 23, 16, 27, -18, 75, 54, -128, 98, 93, -16, -36, -38, -60, -65, 54, 57, 26, 22, -76, -128, 32, 37, 76, -13, -128, 88, 15, -39, 80, 54, -57, -92, 103, 107, -128, 2, 26, -58, 49, 127, -88, -123, 127, 27, -52, 0, -28, 26, 32, 69, 10, 13, 98, -109, 29, 107, -50, -128, -49, 59, 102, 6, -60, 27, -22, 13, -21, 13, 91, -1, -31, 32, 31, -109, 92, 114, -128, 52, -55, -74, 91, -34, 96, -28, -93, 117, -58, -113, 127, 3, -81, 66, 42, 10, -124, 70, -5, -113, 54, 95, 18, -7, -48, -85, 102, 10, -106, -5, 73, 13, 33, 113, -29, -47, -52, 96, 16, -102, 127, -37, -44, 23, 58, -32, 44, 92, -128, -75, 8, 71, 127, 0, -113, -50, 113, 103, -92, -22, 66, -48, -17, -75, -49, -16, 52, 32, -119, -64, 127, -32, -73, 74, 1, 121, 7, -128, 76, 47, -92, 54, -55, -71, 87, 6, 10, 1, -23, 127, -52, -92, 122, 106, -32, -128, -26, 50, 81, -31, -44, 34, -32, 15, 55, -42, -37, -68, 47, 7, -128, 6, 73, -36, 49, 109, -59, 28, 78, -96, -28, 55, -31, -107, 47, -33, -33, -31, 47, 16, -31, -7, -85, -12, 39, -15, 122, 117, -116, -7, -10, -53, -52, 73, 44, -33, -15, 34, -13, -73, -6, -11, 12, -28, 79, 8, -31, 12, 8, -13, 60, -52, 7, -52, -33, 16, -36, 76, -22, 65, 16, -1, -17, -2, 38, 55, -69, 54, 60, -52, -48, 64, 69, -66, -128, 34, -26, 24, -2, 13, 0, -76, 13, 18, 47, 93, -13, -21, 127, -45, -128, 21, 127, -37, -12, -7, 49, 71, -128, -2, 50, -2, 29, -13, -37, 88, -31, -31, 81, -23, 118, 31, -112, -66, 81, 70, -23, 36, 37, -60, -128, 103, 73, -27, -112, -53, 15, -28, 28, 42, 80, 27, 6, 80, -16, -42, -27, -16, 59, 1, -50, 1, -80, -128, 127, -50, -29, 78, 15, -1, -128, 91, 49, -33, 29, -29, -121, 55, 75, -122, -78, 21, 103, 63, -96, -27, 52, 52, 91, -85, -59, 91, -71, 34, 93, -128, 34, 31, -47, 42, -128, 29, 80, -45, -13, -23, -44, 64, 1, -127, 127, 36, -128, 65, -33, -32, 127, -32, 8, 44, -64, -59, -21, 81, -55, -64, -22, -8, 127, 64, -128, -96, 127, 93, -6, -87, -66, 127, 92, -96, -128, 96, 127, -128, -34, -29, 27, 64, -31, 27, -26, -65, 127, 88, -128, -27, 54, -26, 97, -17, 68, 66, -128, 16, 23, 44, 45, -73, 13, 22, -128, 55, 88, -128, -48, 60, 11, 95, 74, -28, -76, 78, 60, -128, 29, 76, -44, 32, 18, 21, 3, -88, -45, 76, -122, 8, 92, -44, -73, -28, 8, -13, -3, -58, 49, 59, -48, 29, 123, -6, -7, -128, -42, 85, -63, -42, 3, 91, 107, -5, -65, -3, -42, -80, 81, 32, -102, 38, 18, 21, -42, 59, -24, -34, 127, -27, 12, -90, -112, 127, 102, -128, 69, 28, -57, -23, -2, 81, 32, -74, -36, 18, -68, 98, 53, -15, -66, 2, -7, -15, -5, -17, 11, -18, 100, -68, 3, 81, -128, 48, 53, -128, 96, 70, -121, 6, 55, 32, -108, -22, -10, 52, -54, -47, 119, 29, -74, -85, 65, 95, 13, 26, -102, -87, 58, 7, 42, 10, 101, 49, -128, 18, 90, -73, -64, 127, 47, -38, 22, -128, -8, 22, 54, 48, -54, -1, -55, 66, 27, -22, -13, -70, 34, 58, -43, 42, 34, -32, 42, -37, -118, 102, 96, -58, -128, -85, 127, 97, -128, 3, 121, -50, -2, -1, -117, -6, 5, 24, 7, 64, -28, 2, 127, -24, -114, -28, 48, 100, 73, -108, -74, 127, -36, -114, 127, -7, -64, 65, 121, -60, -128, 106, 107, -128, -32, 21, 5, 88, -5, 1, -43, 16, -24, 95, 127, -128, -112, 38, 127, 75, -119, 42, 53, -103, -81, 43, 86, -31, 76, 7, -42, -60, -22, 96, -48, 58, 64, -52, -28, -55, -17, 103, 74, -75, 21, 66, -47, 24, 54, 69, -96, -10, 79, -10, -128, 28, 0, -28, -11, -57, 8, 123, -3, -43, 18, 0, -15, 96, 80, -97, 8, 52, -128, -50, 127, -33, -13, -49, -124, 93, 29, -22, 49, -23, -2, 79, 121, -33, -128, -27, 107, -2, 43, 70, -55, -114, -65, 127, -48, -119, 101, -28, 112, 44, -113, 88, 60, -128, -118, 127, 70, -119, -64, -13, 54, 45, 32, -22, 43, 42, -81, -26, -74, 12, 53, 44, 13, -42, -6, -2, -3, -127, 18, 74, -49, -102, 27, 43, -39, -121, 43, 58, -63, 93, -6, -16, -36, -88, 10, 37, -34, 107, 127, -128, -55, 64, -44, -10, 31, 124, 122, -128, -116, 127, 81, -28, -128, -3, 44, 8, 8, -109, -44, -1, -3, 124, 96, -73, -128, -27, 127, -42, -119, 127, 12, -39, 0, 0, 85, 0, -52, 70, 28, -31, 45, -2, -29, 96, 108, -15, -70, -18, 71, -1, -52, -109, 7, 74, -5, -17, 13, -38, -27, 50, -106, 36, -18, -73, 5, 73, 63, -76, -53, 123, 24, -59, 88, -15, -128, 79, 0, -13, 28, -63, 33, -11, 3, 127, 29, -128, 23, 76, -17, -34, -27, 95, -49, -16, -10, -11, 23, 59, 45, -60, -12, 102, 33, -124, -48, 112, -97, -16, 64, -57, 54, 47, -79, -118, 91, -17, -97, 63, 68, 17, -2, -128, -1, -22, 22, 101, -87, 36, -12, -128, 6, 127, -85, -93, 76, 65, -33, 10, 15, 39, 111, -128, -24, 59, -45, 12, 50, 11, -122, 5, 81, -114, 68, 28, -107, 79, -23, 24, 65, -28, 5, 42, -55, -26, -81, 50, 6, -87, 29, 33, 113, -76, -38, 54, 12, -96, -66, 97, 95, -52, -95, 42, 49, -76, 81, 79, -48, 47, -70, -98, 70, -33, -24, 23, 117, 5, 44, -73, -27, 43, -6, 52, -1, -57, -27, 42, 23, 18, 109, -79, -1, 127, -66, -128, -42, 45, 127, 43, -106, -78, 127, 80, -128, -79, 127, 109, -106, -16, 65, 1, -5, -118, -58, 23, 1, 26, 12, 13, -128, -11, 127, 2, -58, -68, 71, 11, -52, 23, -78, 38, 79, -128, -12, 127, -78, -75, 109, 13, 42, -22, -97, 68, 34, -21, -106, -76, 57, -59, -50, 106, 63, -114, -5, 33, 13, 12, 57, 97, -13, -31, -39, -69, 53, -86, -69, 5, 34, -11, 52, 47, -3, -54, -18, 81, -65, 71, -45, 0, 127, -128, -70, 74, -44, 36, 57, -38, -128, 1, 88, 55, -59, -88, 37, 2, 2, 85, -21, -128, -42, 60, 87, 66, -44, 55, -47, -59, 98, -60, -69, 91, 6, -3, -52, 12, 21, -128, 5, 71, 6, -103, 12, -22, 5, 1, 10, -1, -49, 21, 37, 22, 29, 95, 57, -23, -26, -106, -31, 81, 8, 32, -24, -97, 59, 121, -114, -52, 21, 91, -31, 37, 121, -49, -128, -8, 127, -34, -39, -98, 15, 127, -108, -128, 113, -17, 43, 33, -92, -18, 127, 53, -16, -96, 7, 31, -128, 93, 95, -128, -13, 114, -113, -28, 96, -75, -69, 90, 87, 3, -39, -73, 22, -117, -5, 81, -103, 6, 127, -59, -44, 76, -121, -10, -6, 87, -29, -108, 127, 73, -93, -63, 50, 11, -124, -8, 127, -57, -119, 106, 0, -128, 60, 31, -47, 3, 124, -15, -18, 54, -23, -75, -2, -93, -75, 127, 109, -128, -118, 127, -33, -11, 47, -118, 29, 100, 7, -32, -93, 111, 18, -63, -49, 93, 106, -128, -79, 93, 73, -128, 11, 79, -8, -42, -1, 69, -73, -7, -37, 6, 80, -42, -36, 127, -23, -37, 39, 36, -102, -17, 116, -50, -114, 96, 8, 21, -64, -37, 85, 18, -12, -101, -12, 6, 53, -45, -79, 127, 58, -128, 7, 5, 6, 86, 93, -27, -128, 18, 38, -32, -29, 0, 113, -7, -102, 7, 43, 8, 85, 97, -128, -44, 26, 16, 76, 28, -59, -11, 31, -128, 55, -11, -100, 31, 106, -37, 34, -54, 11, 44, -57, -48, 75, 23, -47, 109, -18, -12, -58, -49, 116, -27, 18, 90, -18, -78, 3, -28, -59, 45, 31, -54, 44, 68, -53, -26, -86, 11, 95, 42, 5, 5, -15, -96, -86, -10, 22, 71, 90, -88, 11, 5, -63, 22, -39, -31, -24, -24, 116, 29, -10, -49, 26, 23, -118, 3, 127, -88, -12, 69, 6, -16, -58, 42, -102, 31, 127, -112, -71, 98, 18, -92, -29, 7, -57, 107, 91, -114, -97, 70, 114, 6, -8, -34, -106, 69, 103, -128, 33, 58, -48, 29, -95, -55, 85, -18, 111, 10, -78, 27, -24, -28, 114, 58, -71, 43, -11, -96, -38, 66, 90, 42, -103, -33, 37, -8, 2, -13, 57, -12, 74, -21, 26, 117, -109, -87, 127, -29, -43, 36, 7, 66, -22, -55, -8, 124, -64, 7, -2, -71, 43, 97, 107, -91, -116, 7, 97, 2, -36, -42, 39, 6, -32, 36, 127, -6, -79, 85, -5, 10, 69, -7, -100, -66, -32, 88, 5, -65, 64, 12, -2, 76, -66, -11, 17, -3, 111, 63, -11, -124, 71, -1, -108, 127, -15, 15, -28, -43, 68, -3, -43, 2, 17, 33, 50, -45, -75, 90, 23, -42, -74, -95, 66, 34, 7, 32, 18, -57, -17, 38, -5, 127, -12, -124, 127, 22, -128, 127, 113, -102, -54, -44, -66, 127, 103, -45, -81, -87, 95, -48, 48, 127, -128, -60, 32, 31, 86, 1, -55, 34, 10, -73, 6, 27, -39, -44, -86, 36, 49, -108, -11, 3, 23, 33, 113, -47, -127, 59, 42, 81, -17, -86, 81, 3, -11, -81, -76, 106, 97, 0, -55, -6, -21, -17, 31, 114, 49, -86, -24, -33, 24, -91, 0, 18, -23, 81, -16, -12, 92, 12, -108, -42, -18, -15, 127, 81, -128, 50, -8, 0, 18, -34, -37, 8, 80, -37, -52, 16, -70, -47, 13, -33, 38, 127, -66, 5, 13, -32, -17, -28, 11, 49, 42, -58, 23, 3, -92, -71, 66, 74, 63, -111, -75, 55, 98, -45, 48, 12, 1, -53, -1, -13, -55, 27, -39, 95, -17, 3, 29, -27, 112, 10, -128, 38, 3, -100, 54, 90, -57, 91, -33, 36, 117, -128, -85, 78, 29, -66, -43, 65, 55, 69, -1, -10, -101, 8, 52, -88, -15, 93, 39, -103, -29, 106, -117, -15, 127, -92, -103, -28, 28, 59, -23, -8, 117, 5, 36, -49, -29, 127, -36, 15, 22, -128, 36, 100, -6, -108, -102, 26, 15, -50, 101, 122, -128, 36, 96, -128, -23, 127, -73, -24, 29, -66, 101, 96, -71, -58, 76, 53, -128, -73, 123, -95, -28, 109, 36, -48, -128, -32, 127, -3, -116, 79, -16, -60, 65, 88, -87, 10, 58, -108, -23, -65, 44, 23, 59, -58, -3, 108, 26, -128, -103, 127, -57, 2, 92, -128, -12, 127, -33, -53, -5, 68, -24, -12, 127, 7, -102, -57, 71, -32, 31, -2, -66, 44, 50, -37, 16, 16, 101, 11, -114, 127, -23, -121, 127, 76, -100, -86, 75, 64, -24, 37, -64, 1, 12, -58, 42, 88, -1, 60, 44, -128, -76, 127, 10, -76, 107, -2, -70, 7, 39, -28, -34, -119, 69, 37, -8, -60, -13, 34, 12, 95, 21, -60, -80, -100, 76, 74, -42, -102, 21, 33, -71, 79, -8, -7, -6, -37, 17, 98, 107, -128, -44, 101, -57, -27, 127, 68, -121, -42, -31, 112, 22, -128, 80, 118, -111, -37, 57, 44, -3, -118, -55, 121, 75, -97, -65, -66, 60, 68, 0, -29, -15, -54, -86, 124, 31, 33, -3, -36, -38, -5, 44, -5, 5, -71, -2, -73, 87, 2, 1, 49, -85, -64, 33, 23, 36, -85, -11, 68, 15, -23, -97, 31, 97, -45, -63, 127, 123, -100, -52, -29, -52, 22, -5, -34, 127, 106, -128, 13, 127, 16, -128, -58, -13, 78, 100, -128, -118, 118, 69, 11, 42, -37, -128, 3, 113, -58, -32, 101, 37, 27, 16, -22, -127, -124, 127, 117, -70, -13, -44, -45, 33, 17, -128, -116, 127, -27, -114, 127, 37, -54, -16, -33, -60, 26, 86, 0, -43, -124, -13, 47, -64, 33, 33, -12, 44, -24, -11, 26, -28, 127, -50, -128, 127, -10, -111, 122, -6, -66, 70, -85, -69, 64, 57, 3, -108, 27, 54, -128, 102, -10, -59, 5, 33, 111, -37, -98, -50, 127, 43, -112, 90, 23, -86, 59, 44, -37, -13, -76, -53, 66, 13, 10, -66, -39, 47, 23, -44, -52, 102, 5, -53, 127, -39, -29, 90, -48, 6, 5, -78, -63, -53, 21, 127, -3, -117, 69, -10, 45, 107, -96, -63, 5, -52, 45, 78, -36, -107, -100, 108, 112, -128, 42, 91, -128, 1, 43, -128, 42, 59, -32, 95, -44, -22, 34, -16, 16, -95, -128, 117, 22, -39, 0, 38, 60, -128, 3, 54, -79, 39, -33, -85, -53, 38, 15, 7, -7, 69, 11, 1, -45, -128, 127, 86, -23, -33, -45, 44, -118, 7, 109, -64, -43, -24, 27, 28, 21, 1, -49, -6, 52, 93, 23, -32, -64, 70, 112, -106, -34, 7, -70, 96, 6, -128, 66, 12, 21, -10, -97, 101, 112, -17, -128, -45, -11, 64, 97, -42, 33, 13, -58, -91, -5, -3, 52, 64, -128, 49, -8, 29, 5, -48, 96, 22, -34, -55, 90, -45, -34, -16, -79, 107, 127, -107, 6, 97, -52, -71, -59, 33, -26, -90, -44, 127, 21, -22, 10, -57, -3, 31, -58, 31, -48, 68, 23, -52, 1, -43, 100, 79, -114, 7, 8, -88, -44, 48, 39, -65, -12, 127, 81, -70, -128, 90, 39, -75, 54, -85, -81, 60, 127, -27, 42, 66, -128, -48, 44, 42, 42, -52, -12, 127, -97, 26, 28, -111, 44, 79, -39, 0, 59, -71, -38, 109, 127, -28, -128, 52, 86, -114, 81, 12, -90, 93, 91, -90, 12, -63, 3, 23, -85, -17, 13, 37, -43, 53, 64, -29, -64, 53, 107, -55, -28, -112, -63, 127, 34, -73, -10, -12, 31, 17, 8, 78, 80, -76, -128, 127, 57, -128, -5, 127, -58, -21, 11, -49, 0, 87, 54, -95, -36, 45, -100, -54, 112, -26, -119, 10, 98, -15, -33, -66, 33, 111, -21, -59, -102, 70, 12, -33, 52, -23, -37, -121, 5, -15, 26, -23, -65, 113, 57, 31, -37, -128, 28, 85, -5, 23, 63, -85, -108, 59, 24, 63, -27, -111, 32, 68, -69, -90, 87, 12, -81, 57, 69, 36, 8, -101, 44, 78, -17, -73, -2, -26, -31, -26, 88, -68, 27, 121, -121, -90, 24, 123, -78, 28, -17, -13, 65, -57, -116, -2, 127, -85, 22, 24, 6, 0, -44, 42, -54, -11, -21, 118, 75, -85, -86, 27, 65, -88, -6, 127, -63, -12, 68, -90, 5, -86, -52, 80, 33, -52, 45, -8, -85, 37, 45, -88, -96, 31, 127, -36, -31, 98, -96, -70, 45, 16, -71, -43, 127, 55, -100, -49, 95, -18, 57, 47, -73, -23, 127, 96, -109, 7, -28, -128, 76, 26, -50, 96, 27, -97, -55, 48, 11, 26, 92, 27, -128, 49, 119, -58, -69, -117, 90, 127, -128, -28, 49, -43, 80, -7, -63, 23, 10, 85, -1, 36, 79, -64, -44, -26, 36, 12, -8, -128, -74, 114, 76, -95, -32, 80, -101, -93, 127, 123, -128, 26, 60, -92, -27, -11, 98, 23, -39, 76, 75, -52, -63, 42, -64, -75, 47, 2, -31, 47, 53, 7, 127, -66, -32, 64, 23, 0, -59, -10, -10, -13, -15, -106, 92, 70, -128, -6, 127, -32, -128, 88, -54, 7, 78, -90, -78, -29, 113, 3, -34, 127, 2, -106, 121, -60, -8, 113, -28, -79, -32, 10, -63, -37, 103, -22, 43, 91, -59, -7, -57, -128, 91, 64, 7, -49, 6, 65, -113, -55, -65, 69, 26, -50, 121, -70, -59, 100, -95, -37, 29, 49, 87, -85, 1, -6, -54, 33, -52, -63, 34, 65, -63, -71, 13, -23, 75, -7, -95, 13, -53, 37, 31, -15, 127, -66, -34, 70, -123, 66, 127, -123, -58, 98, 10, -90, -44, 7, -23, -66, -22, 43, 8, 92, 86, -26, 55, -15, -128, -5, 127, -90, 0, 8, -53, 112, -24, -101, 26, 48, 102, -45, -22, 32, -85, 39, -45, 68, -1, -59, 127, -76, -48, 116, 2, -128, -26, 92, 18, -39, -112, 60, 68, 2, 38, -128, 0, 44, -88, 127, 63, -128, -17, 71, 48, 11, 59, -7, -96, -54, -13, 50, 43, 71, -31, -88, 127, 55, -26, -26, -119, 79, -15, -18, 73, -128, 33, 22, -76, 103, -31, -128, 127, 64, -111, 10, -37, 2, 12, 42, 60, -52, 63, 73, 7, -128, 37, 108, -76, 1, -74, 21, 28, -59, -8, -52, 24, -27, 1, -63, -59, 0, -15, 26, 74, 8, -12, 24, -128, -116, 100, 74, -32, -33, 32, 5, -1, 39, -21, -27, 52, 101, -37, -52, 71, 127, 28, -101, -12, 60, 11, 38, 31, -128, -47, 127, 26, -93, 6, 59, -71, -91, 0, 93, -10, 1, -98, 37, 12, -111, 127, 12, -39, 75, -69, 18, 27, -128, -27, 24, 86, 121, -128, -17, 127, -44, -79, 28, 79, -106, -44, 38, -17, 91, -65, -128, 124, 11, 8, 86, -109, -21, -15, -97, 66, 112, -108, -60, 127, -18, -68, 60, -34, 16, 10, -53, 127, 44, -54, 52, -7, -112, -42, 24, -8, 68, 15, -106, 127, -5, 10, -5, 3, -36, -71, 59, -80, 17, 113, 18, -11, -128, -52, 127, 0, -95, 87, -27, 2, 18, -111, 26, 87, -37, 18, -100, -85, 66, -6, -2, 95, -27, 21, 66, -32, -59, -28, 85, 73, 52, -73, -74, 119, 7, -122, -15, 127, -87, -11, 106, -33, -128, -3, 85, 26, -34, -5, 78, -18, -23, -102, -60, 127, 33, -26, -85, 5, 79, -31, -98, 16, -73, 24, 85, -32, -107, -66, 127, -15, 54, 16, -18, 58, -16, -114, -28, -22, 78, -2, -11, 23, -73, -85, 34, 11, -101, 127, -33, 8, 87, -102, -2, 43, -87, -54, 42, -13, 12, -45, 18, 37, 2, -8, -37, 16, 53, 45, -36, -44, -70, 2, 8, -113, -49, 54, 75, -13, -12, 95, -36, 106, -37, -8, 117, -95, -74, 1, 88, 52, -73, -68, -23, -38, 98, 50, -52, -23, -16, -37, -37, -55, -2, -16, 6, 60, -13, 50, 13, -37, -52, 29, 33, -58, 10, -5, 44, 49, -33, -43, -11, -55, -79, -26, 102, -12, -112, 102, -26, 69, 11, -33, -17, 17, 81, -43, -96, -44, 38, 97, 29, -43, -48, -49, -50, -27, 127, -36, -114, 127, 96, 7, -116, -100, 32, -1, 64, 34, 48, 26, -71, -54, 23, 87, 100, -92, -71, 34, 38, 80, 101, -107, -75, 85, 18, -12, 22, -34, -17, 65, -95, -37, 106, -31, -22, 86, -43, -128, 6, 34, 66, 49, -70, 58, 107, -2, -42, -128, -80, 28, 127, -31, -45, 28, 60, 109, -13, -92, -39, 16, -15, 39, 95, 36, -1, -107, 7, -12, -65, 127, -29, -7, -16, -49, 39, -47, 0, 7, -13, 32, 6, -75, 31, 96, -76, -85, 91, -59, 1, 127, -96, -24, 26, -117, 63, 36, -23, 18, 32, 65, -69, 53, 26, -54, -5, -66, -50, 3, 118, 48, 5, -71, 24, 26, -112, -21, 121, 93, -114, -54, 121, -10, 54, -69, -75, 88, -22, 34, 54, 0, -74, -128, 107, -36, 12, 48, -95, 98, 0, 12, -28, -109, -6, 5, 95, -2, -45, 37, -45, 37, 98, 22, 15, -44, 3, -69, -92, 32, -1, -5, 43, 100, -17, 97, 31, -15, -52, -10, 50, -21, -7, -114, -76, -3, 69, 127, -60, 11, -27, -54, 18, 101, -42, -98, 88, 127, -53, -34, -23, -24, 95, -32, 43, 64, -113, -38, 80, 32, -81, -2, 63, -80, 58, 100, -117, -47, 96, 18, 79, 15, -44, -76, -16, 112, -60, 37, 52, -63, -28, 37, 47, 12, -3, -87, -34, -87, 70, -6, -21, -42, 21, 8, -92, 49, 121, -73, -28, 17, 0, 17, 66, -76, -27, 16, 43, 66, -128, -17, 33, 27, -10, -53, 95, -5, 55, 6, -59, 97, 31, -114, 86, 18, -71, -37, 102, 15, -80, 42, 45, 52, 28, -85, 26, -28, -36, 58, -119, 39, -10, -53, 36, -10, 27, 78, -26, -93, -49, 112, 119, -70, -12, 5, 1, -117, 0, 71, -68, -92, -21, 7, 127, 122, -108, -10, -21, -91, 57, 55, -102, 78, -27, -33, 34, 29, 11, 18, 73, -69, -45, 55, 78, -91, -71, 111, -8, -103, 26, 121, -80, -45, 119, -121, -37, 42, 44, 52, -79, -73, -24, 36, -45, -22, -28, 21, -23, 13, 10, 59, 79, -65, -59, 23, 39, 2, -63, -85, -48, -3, 47, 45, 85, -52, -21, 12, 21, 11, -68, -5, -28, -63, 39, 102, 28, -18, -74, 57, -34, -31, 87, 75, -111, -109, 127, 108, 28, -128, -91, 10, 42, 71, 26, -71, 70, -26, -26, 59, 16, -106, -79, 18, 8, 74, 69, 27, -122, -119, 118, 17, -15, 5, -38, 71, 10, 59, 2, -73, -37, 91, 52, -27, -12, -55, 119, 3, -50, 59, 97, -64, -12, -13, -32, 127, 27, -128, 23, 106, -124, -55, -10, 57, 63, -80, -66, 127, -50, -32, 21, -58, 26, 86, 48, -38, 16, -28, -3, 102, 0, -85, -75, 16, 76, 24, -48, -28, 103, -54, -58, 10, 63, 44, 37, -70, 15, -39, -79, -2, 103, 55, -114, 118, -55, -11, 47, -27, 95, 11, -102, -18, -39, 17, -53, 66, 12, -70, 27, -37, 70, 81, -58, -42, 12, 10, 86, -22, -18, 127, -57, -95, 60, 47, -26, 15, 127, -31, -21, 87, -128, -71, 76, 22, -106, 53, 57, -58, -47, 96, 37, -6, -17, 10, 86, -57, 10, -26, -27, -17, -42, 112, 1, -31, 127, -55, -24, 100, -34, -57, 29, 26, 5, -90, -87, 119, -88, 2, 27, -103, 68, 75, 23, 16, -91, -3, -7, 97, 81, -90, 47, 28, -128, -65, 28, 127, -6, -26, 52, 7, -96, -50, 88, -79, 55, -28, -118, 127, 88, -128, 52, -39, -11, 44, -12, 32, -11, -32, -45, -43, -70, 31, -2, -48, 80, -3, -75, -38, 18, 6, -21, 101, 69, 13, 10, -71, 15, 49, -102, -8, -38, -38, 127, 63, -24, -65, -17, 13, -68, -33, -16, 58, -53, 8, 0, -108, 36, 101, -32, 3, 76, -64, -70, 31, -17, 117, 74, -32, -10, -128, -10, 127, -45, -85, 74, -18, -118, 88, 5, 11, 1, 16, 38, -21, -1, 49, 6, 2, -45, 26, -2, -107, -6, 103, 39, -55, 42, 1, -36, 42, 34, 87, -49, 39, -26, 55, -8, -114, 113, 5, 33, 60, 12, -102, -73, 42, 127, 48, 13, -98, -38, 43, -26, 68, 96, -16, 0, -59, 15, 100, -69, 39, -10, -66, 50, -6, -39, 52, 12, 18, 48, -128, -31, 93, -54, 8, 86, 37, 47, -98, -6, -22, -44, 101, 12, -128, -29, 44, -8, 100, 92, -90, -34, -53, 60, -34, -29, -8, 47, -48, 39, 64, -128, 0, 2, -3, 124, 34, 23, -26, -10, -15, -17, -65, -49, 24, -13, 32, 17, -33, -44, -2, -70, -49, -26, 1, 91, 55, -38, -58, 58, -7, -128, -55, 127, -10, -92, 93, 75, -78, -69, 97, 103, -121, -103, 85, 81, 16, -80, -11, 33, -96, 13, -26, 31, 102, -55, -53, 23, 101, 22, -114, -42, 91, -33, -73, -55, 70, 127, -32, -17, -113, -49, 117, -54, -17, 1, -87, 28, 97, 36, -128, -113, 81, 15, 53, -32, 10, -29, 22, 80, 22, -102, -96, 127, 38, -53, 57, -65, -34, 75, -74, 49, -5, -95, 26, 127, 22, -91, 3, 3, -21, 47, 5, 7, 52, -117, -128, 96, 28, 17, -18, -85, 114, 0, 29, -43, -2, 55, -78, -48, -23, 64, -49, -17, 107, -53, -42, -6, 73, -91, 27, 18, -10, 23, -108, 71, 86, -111, -28, -18, 107, 65, -128, 43, -50, -52, 31, -22, 12, 127, 42, -39, -1, 43, -69, -29, 17, 64, 75, 39, -34, -71, -52, 3, -36, 37, 23, 58, 63, -55, 27, -6, -107, -54, 47, 18, 6, 26, -33, 10, -39, 59, -60, -11, 71, -98, -73, 101, 101, -28, -33, -48, -48, -76, 127, 28, -70, -17, -26, 22, 122, -50, 47, -15, -74, 64, 34, -78, -43, 32, 111, 49, -128, 101, 6, -23, -28, -34, 66, -63, -11, 43, 65, 52, -65, 0, 113, -1, -48, -112, 73, 39, -128, 90, 34, -49, -44, -64, 69, 24, -60, 1, -58, 28, 49, -18, -23, 31, 78, -8, -42, -111, -79, 54, 119, -31, 24, 54, -128, 5, 127, -106, -88, 39, 127, 60, -38, -59, -117, 81, -23, 17, 31, -52, 16, 93, 63, -37, -52, 27, 3, -85, 93, 37, -59, 13, 58, -45, -86, 109, 74, 3, -27, -23, -128, 16, 68, 27, -95, -15, 76, -87, -28, 121, -2, -42, 13, 91, 53, -69, -57, -76, 64, -15, -6, -27, 29, 18, -63, 101, -69, -103, 127, 78, -12, -24, -79, -58, 32, 23, -107, -44, 127, -21, 43, -65, -11, 47, -111, 95, -10, 8, 127, 1, -16, -52, -128, 43, 127, -68, -52, -58, 45, 32, 50, 22, -128, 23, -24, 102, -3, -101, 26, 127, 12, 16, 65, -128, -69, 127, 31, -112, -12, 48, -57, 0, 6, -21, 127, 100, -100, -70, -74, -21, 127, 91, -50, 0, -81, -23, 70, -76, 8, 65, -113, -92, 127, -34, -69, 33, -36, 127, 36, -81, 11, 8, 52, -31, -21, 33, -47, -69, -26, 54, 22, 80, -29, -128, 112, 64, -29, -15, -128, 29, 58, -60, 75, -22, -44, -24, 21, 73, -81, 91, 127, -102, -75, 44, 86, -128, -55, 68, -21, 31, 71, -7, -65, -92, 66, 13, -128, 88, 8, -92, 66, 79, 2, -75, 87, 93, -128, -68, 31, 2, -8, 1, 100, 48, -128, 48, 118, -73, -79, -17, 8, 23, -15, 121, 68, -128, 0, 102, 54, -42, 0, -54, -78, 33, 65, -22, -27, 127, 22, -26, -63, 43, 111, 3, -106, 8, 43, -122, -32, 127, -24, -53, -33, 8, 34, 43, -1, 3, -29, -60, 12, -18, 59, 50, -36, 96, -2, -75, 28, 71, -128, -2, 86, 5, -29, 11, 5, -123, -57, 2, 27, 93, 63, -58, 70, 88, -128, -44, 124, -44, 6, 87, -75, -111, 1, 106, -65, 29, -1, -5, 71, -107, -18, 21, -48, -17, 44, 127, -26, -65, 108, -29, 16, -27, -36, 78, -97, -8, 1, -108, -3, 39, -10, 97, 45, -38, 3, 31, -39, 33, 15, -106, -39, 127, 31, -128, 123, 45, -15, -80, -128, 121, 87, -128, -42, 101, -58, 58, 37, -45, 88, -16, -36, 66, -96, -107, 57, 86, 39, -13, -55, -78, 78, 36, -103, -23, 116, -32, 52, 68, -102, 74, -8, -128, -42, 127, 86, -128, 7, -11, 39, 43, 1, -6, -45, 106, 1, -18, 12, -70, -2, 127, -13, -122, 34, 78, -31, 98, 36, -128, 29, 127, -113, -113, 52, 22, 127, 86, -121, -63, 106, 54, -49, -69, -87, 122, -16, -52, 70, 6, 10, 34, -57, 26, 48, -53, -70, -98, 75, 127, -119, -91, 127, -33, -90, 127, -22, -128, 111, 54, -66, 13, -2, -86, 123, 23, 3, -92, 23, 43, -53, 23, -76, 107, 0, 1, 21, -60, 59, -101, -32, -27, 5, 73, -50, 73, 13, -42, 91, -73, -102, 54, 119, 7, -60, 44, 87, -90, -15, 78, -12, -79, -53, 127, -26, -23, 98, 24, -96, 2, 123, -12, -54, -48, -74, 92, 127, -91, -128, 96, 32, -95, -47, 16, 113, 5, 29, 0, -29, 3, -54, -11, 101, 3, 60, 43, -28, -15, -66, 73, 101, 23, -117, -68, 6, 5, -6, -7, 113, 0, -112, 10, 106, -43, -3, 18, 13, -3, 29, 119, -50, -55, 75, 16, -60, -38, -53, -58, 121, -5, -15, 44, -96, -79, -12, 90, 38, -50, -96, 15, 127, -92, -3, 52, -85, -38, 81, 66, -74, -63, 50, 70, 13, -70, -24, 5, -79, -69, 127, -8, -43, 118, -101, -88, 48, 63, 116, 34, -18, 8, -124, 10, -31, -97, 74, 60, -1, -38, -6, 122, 11, 12, 15, -88, -5, 0, 97, 28, -100, 43, 49, 11, -55, -18, 59, -37, -128, 60, 27, 43, 17, -64, 23, -1, -3, -98, -75, 127, -23, -114, 117, 17, 54, -87, -15, 17, -53, 48, 58, 1, -107, -5, 45, 36, -57, -28, 28, -13, 127, 26, -128, 50, -6, 73, -1, -1, 111, -111, -7, 118, -66, -91, 21, 18, 18, -47, 49, 102, -28, -68, -31, 63, 38, -15, -76, -128, -12, 127, -11, -64, 17, 36, 103, -38, 78, 68, -52, -7, 10, -70, -26, -22, 34, -55, 27, 24, -71, 45, 127, 32, -53, -70, -17, 36, -55, -86, 80, 44, -8, 37, -49, 0, -102, -81, 127, 91, -44, -71, -31, 18, -113, -48, 127, 36, -128, 2, 95, -52, -128, 117, 10, -3, -6, 23, 1, -31, -71, -52, 44, 117, -66, 24, 86, -128, -66, 107, -13, 87, -17, -15, 74, -101, -74, 92, 127, -75, -103, 93, 68, -117, 11, -34, -68, 34, -1, 111, 119, -127, 45, -33, 21, 127, -128, -7, 28, -74, 45, 44, -18, 58, -1, 64, 93, -109, -18, 93, 11, 10, -10, -54, 114, -49, -58, 13, -3, 73, 71, 85, -60, -57, -65, 11, 90, -73, -48, 127, -11, -53, 127, -64, -27, 111, -8, -128, 52, -60, -6, 33, -16, -49, 10, 65, -69, -79, 91, 60, -36, -12, 8, 100, 43, -86, -65, -2, 37, 22, -93, 55, 123, -128, -122, 127, -27, 44, 127, -128, -128, 127, 36, -32, 95, -128, -81, 55, -32, 123, 65, -79, -68, -37, 71, -13, 52, 121, -48, -86, 6, 75, -59, -24, 127, -66, 70, 65, -31, 22, -76, -5, 1, -128, 11, 107, -109, 65, -55, -90, 127, 18, -11, -128, 32, 27, -112, 54, 127, -24, -60, -10, -85, 75, 76, -10, -2, -28, -58, 16, 26, -107, 42, 37, -63, 23, -11, 47, 36, -57, 116, -23, 12, 70, -122, 15, 109, -98, 38, 69, -70, -31, -97, 63, -7, 11, 42, -128, 13, 127, 5, -128, -59, 78, 57, -7, 50, 12, 6, 55, -53, -53, -80, 10, 27, -3, -23, 127, 32, -13, 38, -128, -15, 127, -128, 5, 122, -88, 13, -60, -43, 52, -42, 10, 79, -13, -7, -47, -117, 52, 18, 27, -53, -29, 7, -13, 100, -47, -44, 17, -10, 3, 43, 108, -73, -44, 103, -87, -80, 127, 27, 8, -37, 37, 10, -95, 74, 11, 34, 73, 33, -122, -12, 11, 26, 111, -33, -71, 93, 54, -85, -96, -54, 11, 22, 48, 80, 73, -69, -8, 3, 10, -31, -1, 16, -8, 38, 39, -6, -101, 0, 57, -44, 102, 16, -28, 12, 33, -112, -28, 121, -16, -8, 11, -34, 2, -116, -68, 109, -7, 54, -85, -112, 53, 91, 21, 12, -45, -52, 36, 28, 63, 42, -24, -32, 113, -87, 11, 117, -128, -27, 79, 33, -68, -42, 49, -53, 17, 96, 23, -128, 13, 127, -128, -128, 93, 76, 0, -5, -5, 6, 12, -121, -64, 17, 43, -2, -36, 44, -43, 15, -33, 68, 17, -70, 13, -87, 95, -16, 39, 86, -128, 45, 66, -96, 53, -36, -128, 87, 127, -3, -103, 32, -93, 28, 0, -16, -3, -5, -2, -16, -18, -6, 17, 28, -90, -123, 127, -47, -111, 127, 48, -107, 18, -17, 16, 22, -45, 39, -88, -26, 68, 5, -45, 5, 3, -13, -22, -128, 31, -13, 43, -18, -128, 114, 18, -68, 127, -34, -64, 6, -18, 127, 16, -29, -12, -79, 43, -27, -28, 127, 58, 6, -37, -101, 65, -2, -86, 53, 57, -106, 70, 70, -114, 68, -32, -39, -10, -60, 122, 38, -108, 91, 24, -37, 27, 22, 15, 18, -36, -22, -23, -92, 34, -52, 5, 48, -24, -90, -32, 64, 3, -13, 127, 24, 23, -87, 36, -17, -117, 127, 31, -68, -1, 90, 28, -3, -65, -68, 66, -70, -60, 52, 34, -78, 29, 8, 1, -23, -47, -60, 49, 92, -108, 16, 3, -52, 127, -10, -60, 127, 64, -38, -97, -52, 79, 127, -88, -121, 113, -10, 5, 0, 73, 8, -47, 73, 50, -76, 79, -27, -109, 98, 74, -58, -102, 111, 22, -23, 68, -48, -53, 16, -55, 26, 79, -6, -42, 22, 26, -128, 64, 0, -118, 107, 22, -8, -38, 103, 69, -128, -58, 127, 54, -13, -98, 5, 63, -43, -28, -2, -60, 95, 127, -128, -54, 71, 59, -128, -38, 119, -78, -28, 127, -59, 45, -44, -17, -3, -75, 81, 13, 0, 22, 102, 121, -109, -69, 48, 45, 36, -128, 34, 122, -128, -63, 75, 91, -53, -18, 17, 74, 34, -39, 7, 27, -26, -5, -22, -18, 53, 6, -36, 23, 17, -113, 28, -55, 15, 47, -128, 85, 50, 23, -11, -75, -69, 95, -16, -92, 43, 11, 119, 27, -38, -49, -58, -12, -44, 96, 79, -21, -73, -70, 53, -44, 13, 31, -69, 18, -75, 2, 52, 6, 16, -96, -37, 124, 114, -108, 22, -39, -42, 112, 17, -93, -74, -8, 70, 15, -114, 36, 24, 10, -64, -54, 17, -38, 127, 63, -49, -100, -48, 32, 85, 81, -114, 33, 31, -114, -18, 64, 22, 71, -23, -73, 10, 79, 50, -116, -17, -29, 98, 122, -50, -128, -48, 0, 13, 52, 73, 100, -100, 13, -43, -128, 127, 18, 39, -57, -43, -10, 15, 127, -128, -122, 93, 52, 93, -74, -11, 42, -73, 75, 7, 71, 47, -93, 38, 31, -49, -64, 16, -98, -16, -13, -28, 58, 34, -18, 31, -37, 0, 36, -58, 60, 29, -16, 103, -74, -39, 59, -21, 18, 86, -23, -86, 18, -64, -12, 81, -85, -45, 112, -2, 49, 43, -43, -66, -55, 127, 79, -127, -39, -16, 12, 127, -38, -13, 39, -59, -65, -33, -50, 127, 0, -43, 34, 28, 27, -7, -86, -2, -65, -111, 23, 127, 47, -49, -102, 43, 74, -128, -29, 43, 0, 118, -38, 12, 70, 31, -78, 36, -32, -98, 127, -22, 13, -3, -108, 95, -2, 5, 37, -57, 29, 31, -71, -34, 12, 22, -22, -68, 60, 59, -75, 52, -17, -64, 33, 85, -63, -11, 88, -86, 44, 26, -55, 28, 32, -6, -74, -85, 28, 127, -5, -128, 57, -47, 23, 17, 5, -29, -16, 36, 39, 60, -128, 73, -32, -63, 127, -65, -87, 58, 45, 73, 33, -18, -73, -45, 3, 27, 3, -128, 53, 28, -103, 59, 10, -111, 112, -12, -109, 63, 53, -78, -29, 123, 111, -96, -118, 102, 36, -68, -57, 127, -3, -128, 127, 98, -70, -47, 11, -33, -11, 34, -128, -65, 107, 47, -38, -1, 64, 5, -128, -15, 127, -32, -92, 101, 69, -73, 3, -28, 54, 81, -113, 81, 58, 2, 2, -128, 7, 26, 34, -34, -95, 93, 12, -18, -36, -128, 29, 37, 43, 7, -8, -27, 6, 54, -127, -37, 11, 55, 47, 34, -58, -12, 87, 29, -21, -65, 124, -64, -6, 127, -69, -113, 87, -2, -101, 59, 32, 43, 68, -100, -60, 91, 47, 79, -71, -24, 8, -49, 127, 5, -45, 75, -17, -128, -6, -7, -2, 64, -42, -21, 36, 87, 1, -95, 116, 34, -65, -49, 127, -28, -119, 37, 71, 64, 66, -10, -128, 109, 74, -23, -63, -86, 103, -70, -22, 44, -48, -57, 119, 43, -111, -21, -3, 90, -1, 57, 95, -78, -128, 91, 91, -128, -68, 27, 111, 114, -34, -58, 44, -74, -31, -6, 36, 18, -47, -16, 75, 38, -107, 16, -50, 1, -54, -23, 59, -26, 22, -1, 93, -10, -109, 48, 33, -60, 44, -32, -63, 38, 106, -69, -3, 39, -44, 0, 71, 43, -47, -28, -31, -101, 18, -50, -88, 127, 37, -58, -60, -74, 127, -18, -54, 17, 57, -50, -10, 70, -74, 80, -88, -86, 44, 86, 70, -31, -91, 28, 64, -107, 31, 42, -10, 0, 1, 57, -54, -74, 28, 59, -12, -29, 69, 66, -43, -48, -98, -2, 32, 23, 26, -43, 74, 16, 29, -31, -128, -6, 7, 113, 0, 8, -42, 42, -22, -8, 69, -47, -96, -36, 43, 66, 45, 81, -42, -113, 64, 34, 0, 44, 28, 13, -128, -10, 86, -114, -29, 127, -6, -53, 48, 45, -75, 36, 55, -66, 15, -29, 85, 34, -119, 97, 71, -81, 1, -107, 23, 13, -37, 11, -74, 42, 37, -52, 0, -31, 29, 86, 49, -6, 21, -78, -97, 127, 73, -71, -101, -44, 117, -68, 21, -12, -108, 124, 101, -128, 49, 93, -112, 0, -49, 32, -7, -1, 116, -58, -44, -29, -88, 34, 127, 47, -73, -128, 75, 29, -8, -75, 15, 74, -114, 5, 71, -65, -66, 36, -3, -47, -3, -63, -34, 121, 85, -74, -57, 63, 86, -128, -103, 27, 100, -16, 108, -5, -122, 127, 54, -128, -59, 103, 111, -37, -90, 66, -73, 42, 52, -45, -15, -109, 88, 60, -17, -24, 37, -88, -97, 127, -44, -87, 127, 22, -113, 37, 48, -78, -7, -31, -23, 66, -127, -27, 58, -15, -12, 16, -5, 69, -59, 8, -48, -109, 102, 109, 0, -76, 52, 58, -122, -108, 24, 17, 93, 47, -128, 26, 18, -118, 26, 28, -39, 78, 116, -33, 50, -74, -128, 98, 3, 3, 54, -32, 31, 107, 64, -128, -87, 127, -73, -8, 8, -16, -1, -31, 59, 33, 111, 29, -95, -59, 91, 0, -12, 6, 16, 5, -57, 42, -116, 0, 15, -48, 101, 15, -121, 28, 70, -71, -18, 48, -113, 18, 0, -81, -42, 71, 87, 34, -74, -122, 26, 26, 54, 127, 1, -103, 17, -3, -50, 102, -55, -3, 21, 75, -18, -68, 95, -85, -88, 107, -23, -1, 73, -12, 50, 0, -119, 23, 65, -15, 15, 39, -21, 60, -8, -128, 7, 18, 38, 71, 69, -27, -111, -23, 78, 48, 42, -44, -3, 91, 7, -38, -88, -31, -1, -27, 127, -3, -33, 12, 8, 117, 1, -21, 1, -128, 60, -39, -92, 69, 60, -52, 52, 88, -109, -44, 0, 127, 23, -34, 44, -80, -43, 127, 1, -97, 96, -50, -49, 28, -5, -50, 11, 27, 124, -38, -85, 127, -69, -17, 6, 22, 63, 28, -87, 6, -47, -54, 108, 7, -101, -2, 127, -8, -68, -7, 113, -23, -27, 29, 16, 101, -71, -2, 118, -128, 10, 23, -128, 127, 119, -128, -13, 68, -109, 96, 23, -124, 29, -24, 81, 43, -59, 8, 65, 6, -28, -18, 13, 76, -18, -128, 42, 106, -10, -36, -128, 50, -2, -101, 127, 127, -113, -74, 59, -1, -31, 95, 10, -52, 57, -85, -124, 28, 102, 55, 5, -103, -78, 73, -13, 76, 43, -2, 3, -81, -7, 48, -85, -1, 81, 22, -50, -128, 0, 18, 31, 102, -85, -73, 80, 127, -43, -74, 3, -54, 32, 21, 17, 68, 42, -5, -29, -27, 21, 127, 2, -17, 0, -27, -29, -50, 45, -71, 1, -5, -21, 1, 108, 29, -102, 10, 45, 52, 52, 0, -33, 53, -11, -24, -52, -81, 0, 92, 2, -10, 44, 58, -38, -90, 60, 107, -5, -109, 87, -33, -85, 33, -1, -6, 74, 29, -47, 91, 50, -5, -88, -97, 101, -66, -91, 57, 24, 23, 98, -1, 1, -33, -78, 127, -7, -47, 68, 16, 0, -43, -128, -53, 127, -17, -92, 44, 43, 16, -60, -17, 42, 27, 17, -74, -7, 64, -48, -128, -26, 79, 13, 91, -5, -74, 52, 37, -128, -12, 87, 64, -111, -12, 1, -75, 0, 87, 85, 10, -71, -93, 22, 127, 70, -128, -43, 114, -58, -81, 127, 27, -32, -29, -16, 127, 8, 3, 0, -70, -18, -48, 24, 68, -114, 36, 127, -128, -52, 75, 63, -11, -47, -91, 18, 53, -68, 112, -50, -75, -1, 92, 88, -88, 29, 58, -106, -74, 95, 71, -8, -123, -92, 66, -43, -7, 73, -71, 43, 127, -27, -69, 6, -44, 36, -24, 18, 124, -128, 21, 15, -103, 80, 114, -32, -87, 37, 58, -24, -64, 15, -2, 10, -107, -71, -1, 63, 116, -106, -69, 114, 64, -3, -98, 71, 1, -92, 80, -29, -5, 50, -1, 26, 101, -65, -122, 47, 127, 71, -128, -27, 121, 16, -69, 45, -86, -38, 78, 38, -8, -21, -23, -58, 3, 74, -38, 16, 119, -8, -23, -86, 73, 109, -91, -1, -92, 5, -6, 91, 45, -128, 50, 10, 63, 96, 3, -32, -121, -29, 36, 66, -106, 23, 127, -128, -78, -31, 106, -11, -10, 49, -65, 50, 1, 60, -1, -57, 36, 21, 0, 95, 3, 0, 73, 57, -81, -34, 54, -5, -98, -42, 92, -5, -49, 78, 60, -12, 13, -32, 5, 127, -33, -70, -5, 18, -39, 1, 98, -55, -6, 66, 5, -12, -112, -34, 74, 3, -102, -3, 28, -23, 68, 69, -59, 6, -49, 52, -37, -2, -10, -1, 106, -12, -85, -36, 36, 53, 79, 81, -12, -106, 34, 43, -108, 102, 122, -63, -69, -95, -36, 127, -2, 0, 7, -11, -23, -7, 7, -29, -44, 27, -63, 92, -16, -128, 127, -31, -93, 73, 81, 28, -63, -58, -63, 48, 11, -74, 36, -47, 6, 116, 37, -6, -60, -68, 31, -53, -44, 49, 92, 23, 26, 17, -80, 39, 38, -88, -107, -21, 127, 112, -128, -13, 85, -54, -17, 107, 3, -32, 48, -128, -32, 118, 24, -127, -86, 88, -1, -15, 87, 58, -1, -64, -34, -29, 6, 12, 57, 15, -37, 43, -6, -10, -23, 87, 68, -73, 15, -39, -53, 74, -8, -118, 57, 47, -65, 88, 81, -100, 60, -7, -128, 92, 106, -75, 29, -86, -8, 55, -36, -58, -54, 127, 43, -111, 60, -23, 34, 26, -33, -28, -54, 127, -31, -27, 3, -44, 48, -69, 74, 58, -68, 75, -47, -76, 50, -6, 33, -10, 59, 127, -123, -5, 87, -47, 39, -69, -17, 44, -12, -81, 26, 88, -127, -122, 92, 54, -29, -76, 36, 10, 11, -39, -69, 127, -2, -68, 124, 0, -91, 6, -2, 6, -29, -52, 10, 21, 75, -58, 97, 31, -112, 113, -34, -17, -38, -79, 68, 107, -43, 52, 87, -42, -128, -97, 127, 7, -29, 54, 59, -128, -73, 88, 52, 11, -13, 32, 22, -128, 24, 88, -74, -96, 43, 88, 0, -47, -1, -111, -54, 6, -24, 60, -23, -11, 79, 74, -13, -128, 15, 76, -80, 57, 113, -37, -108, -15, 47, -74, 43, 39, -122, 0, 123, 57, -109, 6, 63, -100, 96, -44, -60, 37, 27, 48, -5, -69, 7, 10, -17, 127, 34, -111, 18, 33, -97, -54, 27, 127, -13, 38, -27, -86, 8, 127, -57, -66, 101, 13, -10, -21, 22, -103, 47, 17, -23, 8, -17, -45, 31, 119, -107, -47, 38, 92, 100, -108, 26, -49, -95, 42, 127, -7, -73, 0, -17, 66, 48, 50, -95, -75, 59, 106, -44, -91, 8, -36, 97, 107, -116, -48, 90, -22, 16, 76, 58, -79, 21, 53, -119, 63, 64, -128, -58, 22, 49, 34, 57, -76, -47, 127, -38, -16, 66, -31, -118, -78, 127, 93, -23, -17, 32, -128, 10, 18, -22, 37, -28, -10, -63, 70, 0, 32, -88, -28, 23, -6, -22, 92, 50, -102, 54, 63, -128, -12, 63, -70, 43, -6, -93, 49, 127, 54, -114, -13, -37, -85, 32, 111, 17, -60, 2, -97, 1, 92, -10, -5, -113, 16, 53, -29, -96, -26, 65, -27, -71, -27, 100, 87, -88, -3, -38, -50, 81, 43, -98, -91, -7, 127, -32, 39, 37, 1, -65, -96, 127, 100, 11, -16, -59, -48, 3, -124, -43, 79, 24, 0, 21, -52, -28, -13, -45, 109, 68, -128, 37, 1, -74, 127, 81, -118, 5, -12, 80, 54, -128, 29, 38, -75, 44, 10, -93, 58, 63, -1, -57, -24, 27, 127, 36, -31, -73, 43, 44, 5, 37, -128, 38, 98, -23, -54, -128, 13, 127, -81, -88, 127, 60, -78, -66, -27, 127, -45, 0, -2, -16, 76, -79, 0, 17, 7, -60, -22, 18, 12, -26, -98, 97, -16, -128, 103, 106, -128, -79, 97, -16, -29, 64, 75, 24, -33, -128, 42, -49, 68, -12, -36, 116, -65

);
 
    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project
 
    constant SCENARIO_ADDRESS : integer := 0;    -- This value may arbitrarily change
 
    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
 
                o_done : out std_logic;
 
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;
 
begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
 
                o_done => tb_done,
 
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );
 
    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;
 
    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
 
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
 
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;
 
        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
 
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;
 
        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';
 
        -- Wait some time for the component to reset...
        wait for 50 ns;
 
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
 
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock
 
 
        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
 
        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
 
        wait until falling_edge(tb_clk);
 
        memory_control <= '1';  -- Memory controlled by the component
 
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
 
        tb_start <= '1';
 
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        wait for 5 ns;
 
        tb_start <= '0';
 
        wait;
 
    end process;
 
    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin
 
        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';
 
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
 
        wait until rising_edge(tb_start);
 
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;
 
        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(signed(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;
 
        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);
 
        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;
 
end architecture;

