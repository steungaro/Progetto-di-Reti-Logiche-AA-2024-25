--Testbench created to:
-- -test the component under different input scenarios
-- -test that the result is truncated correctly
-- -test that the component works correctly even after recieving the reset signal mid-elaboration
-- -test both the 3rd order filter and 5th order filter
-- -ensure that the 3rd order filter works correctly even when the first and last coefficients aren't set to zero
-- -ensure that the component can start the conversion again without needing the the reset signal
--This is done by using the example data from ESEMPIO 3 and ESEMPIO 4, which are tested in succession
 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
 
entity tb2425 is
end tb2425;
 
architecture project_tb_arch of tb2425 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
 
    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");
 
    -- Scenario 1
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 12000;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;
    
    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                               -- S
                                                      0, -1, 8, 0, -8, 1, 0, 1, -9, 45, 0, -45, 9, -1           -- C1-C14
                                                      );
    signal scenario_input : scenario_type := (50, 99, 107, 1, -120, 36, 3, 28, 6, -109, 81, -109, 60, -29, 65, 65, -107, -117, -19, 48, -95, -38, 86, 80, 31, -29, 29, 1, 87, -122, -105, 42, -36, -80, 0, 79, -117, -37, -79, -109, 120, 35, 62, 70, -71, -36, 10, -65, -71, -7, 44, -47, 91, -86, -19, 118, -75, -60, -114, 26, -125, -97, -8, -124, -73, 52, 123, 88, -39, 122, -27, 0, 47, 66, -35, 91, 107, 103, -80, 127, 88, -50, 73, 126, 121, -128, 103, 92, 59, -107, -71, 74, 8, -115, -96, 13, -116, -59, -99, 93, -46, 82, 3, -83, 101, 30, 110, 41, 88, -101, -64, 115, 45, 117, 58, -25, -57, -52, 108, 118, -24, 29, -106, 3, 52, 84, -53, -82, -75, 27, -41, 15, -122, 93, 77, 106, -10, -73, 37, 20, 35, 67, 12, 51, -39, -83, 93, -79, 111, -68, -94, 6, -55, 91, -126, 67, -14, -72, -7, -62, 0, -54, -36, 108, 54, 121, 64, 37, -13, 58, 96, 36, -32, -91, 121, 102, -89, -32, 125, 114, 71, 72, 29, 89, -47, 79, -20, 20, 74, 1, 101, -127, 15, 13, -88, -107, -59, -57, -84, -1, 21, 8, -37, 118, 26, 122, 69, 6, 111, 74, 32, 73, 34, -56, -53, 82, 72, -87, 39, -119, -23, 94, 93, -95, 69, 118, -72, -45, -64, -99, 118, -39, -78, 83, 75, -27, -104, -43, 85, 124, -57, -43, 76, -32, 5, -53, 9, -72, -52, -86, -9, 54, -97, -46, -13, 21, -67, -127, 3, 86, 6, -94, -31, -10, 120, -52, 70, -68, -116, 114, -27, -113, 14, -45, -82, 116, 15, 111, -110, 76, -98, -87, 109, -67, 86, 86, 8, 13, -10, -24, -48, -110, -106, 8, 109, 30, -43, 108, -90, 38, -53, -101, -37, -15, 6, 54, 0, 108, -43, -102, -3, 116, 103, 116, 48, 86, 122, 119, -104, -6, 67, 95, -50, -115, -62, 73, -101, 4, 127, 13, -25, 71, -90, -83, -5, 122, -22, -112, -117, -11, 86, 59, 46, 10, 123, 47, -48, 11, 5, 40, -4, -6, 3, 104, 105, 39, -62, 27, -64, 65, -67, 0, -123, 86, 57, 13, -1, -27, -43, -16, -70, 63, 127, 107, -111, 59, -57, 28, 0, -81, 0, -75, -54, 28, -58, -36, -78, -94, 21, -13, -26, 3, 11, -20, 126, 127, 47, -5, -67, -101, -27, -57, -96, 56, -93, 51, 21, 105, -107, -31, -72, -66, -118, 96, -8, -47, 114, 116, 70, -15, -54, -97, -82, 115, -38, -16, 25, -67, 95, -38, -54, 89, -121, -61, -87, -9, -107, 66, -6, 77, 84, 42, -108, -27, 65, -121, 123, 36, -71, 69, 9, -51, -24, -116, 47, 108, 72, -107, 62, 120, 13, 125, -77, -80, 120, 116, -41, 66, 60, 61, 65, 0, 113, -2, 65, 24, 116, 48, 105, -3, -53, -68, 72, 67, -106, 101, -113, 74, -122, 14, 46, 115, 48, -80, -39, 80, -126, -127, -21, 58, 97, 102, -107, -12, -92, -21, 35, 9, -3, 53, -17, 13, -92, -42, -118, -32, 117, 12, 57, -122, 94, -20, 116, 39, 37, 69, -126, 83, -71, 51, 4, 81, 121, -48, -43, -5, -65, -9, 41, 112, -41, -126, 43, -2, -115, -124, 121, 101, 63, -82, -12, -88, 13, -98, 108, 110, 66, -4, -15, 74, -14, -45, -67, -67, 124, 98, 14, -92, 84, 93, -71, -123, 62, 40, 100, -52, -50, -74, 113, 42, 42, -23, -3, 45, 94, 65, 17, 64, 84, 79, 68, 99, 110, 98, 108, 73, -52, 17, -93, -61, 123, 11, -49, -76, -78, 117, -51, -126, -118, -36, -24, 92, 117, -3, 105, 98, 62, -43, 56, -67, 16, 27, -37, -128, 15, -16, 34, -40, 39, -25, 27, -74, 84, 105, 24, 25, 33, -81, 96, -36, -23, 48, 55, -49, 53, 78, -107, 110, -35, -97, -63, -35, 65, 42, -118, -96, 12, 48, 114, 76, -44, 30, -22, 53, -73, 14, -33, -97, 50, 31, -1, -30, -25, -11, 0, 104, -102, 111, 95, -1, -78, 24, -109, 60, -22, 11, 23, 71, -42, -2, -84, -73, 90, 74, 21, 31, -84, -84, 24, 105, -6, -58, 31, -80, 15, 124, -109, 15, 83, -18, 109, 64, 17, 45, 109, -8, 108, 85, 108, 84, -90, -41, -83, 78, -19, -110, 23, 61, -19, 110, 36, 63, -13, 18, -105, 3, -91, 9, 59, 8, 6, 110, -114, -39, -31, -71, -10, 34, -37, -11, -6, 83, -10, 107, 113, 52, -3, 15, 27, 0, 74, 45, -89, 34, -106, -102, -66, 51, -63, 76, -126, -19, -47, -17, -112, -29, -109, 35, -9, -59, -25, -97, -104, -54, 2, 107, -89, -81, -115, 111, 127, 55, -5, -97, 100, -81, -125, 109, 48, -41, -118, 41, -128, -126, 71, 37, 3, -45, 5, 94, 65, 63, 95, 19, -42, 82, 23, 97, 75, 54, -14, -25, 117, -38, 83, 77, 97, -95, -71, -26, -120, 108, 3, -78, 115, 33, -7, -20, 13, 94, -102, 65, -42, 126, 115, -81, 2, 36, -20, -103, -41, 77, 12, 121, 33, 111, 20, 6, 6, -124, -77, -44, 117, -24, -22, 94, 10, -109, 12, 5, -43, 0, -120, 61, -110, 105, -87, 22, 5, -54, 94, 78, -108, -122, -11, 51, 45, 51, 45, 113, -14, 12, -7, -109, -5, -90, -81, -121, 13, -44, -65, -65, 60, -110, -89, -20, 57, -4, -21, -24, -54, -65, -126, 110, -39, 14, 43, 20, 19, 10, 64, -45, 50, 109, 35, -101, 106, -83, -94, -110, -64, -68, -6, 88, -96, 48, 93, 21, -88, -42, -1, -64, 41, -127, 7, -24, 58, 7, -38, -34, 27, 42, 59, -50, -2, 69, -124, -29, 20, -55, 23, 41, 82, -21, 53, -51, -48, 125, -39, 19, 41, 98, -111, 8, -117, -96, 74, 41, 60, -65, 38, 31, 3, -18, 26, -68, 108, 85, -56, -2, 42, 100, -113, 114, 85, -16, -55, 77, -65, 46, -107, 76, -37, 36, -10, -22, 44, -39, -88, 73, -120, -42, 89, -20, 102, -96, -65, 53, -58, 106, 47, -60, 100, -27, -15, -15, 16, -98, 38, -64, -47, -12, 111, 17, -46, 91, -44, -68, 21, 4, -115, -108, -55, -62, 103, 78, 18, -115, -108, 105, -19, -14, 81, -125, 115, -123, -108, -28, -20, -125, -32, 62, 77, -44, 14, -46, -61, -8, -52, -10, -42, 54, -86, 49, -18, 97, -77, -113, -4, 105, -77, -112, -125, -15, -8, 48, 23, -84, 2, 22, 112, -32, 118, -24, -73, 28, 69, -126, 86, -115, -76, -104, 111, 36, 60, 59, 41, -33, -83, 45, 56, -100, -31, 119, 92, 112, -18, -78, -35, -113, 2, -128, 88, -23, 122, 110, 26, -57, 35, 29, -95, 48, -51, 101, -113, -23, -46, 109, -118, -86, 64, 32, 61, 90, 126, -37, 48, -21, -13, 107, -107, 37, -5, 56, 91, 18, 87, -72, 85, 36, 76, 81, 25, 40, -114, 62, 19, 39, 24, -26, -112, -5, -73, 10, 75, 31, 108, -52, 50, 44, 69, -18, 113, -128, -11, -98, -15, 49, 85, -103, 84, -60, 30, -61, 40, 77, 40, 76, -81, 93, -17, 67, -48, -30, -107, -8, 104, -77, -85, -10, -37, 24, 69, 123, 85, 74, 34, -85, -113, 79, 123, -111, 51, 55, -34, -99, 117, -14, -4, 70, 13, -39, -41, -60, -40, -99, 76, -49, -9, -110, 53, 118, 2, 65, -88, -77, -13, 126, -121, 120, 66, 67, 19, 93, -114, 99, -120, -84, -96, 99, 72, -101, -20, 94, 24, -111, -36, 4, 55, -96, 121, -108, -60, -121, 43, -106, -96, 103, -97, -127, -14, 94, 102, -6, 79, 91, -30, -45, -127, 84, -68, -57, -88, 125, -127, 59, 34, 39, 87, 71, -30, -32, 66, -102, 79, -51, -126, 2, -5, -123, 47, 71, -105, 21, -103, 67, 97, -71, 22, -107, 96, -44, 30, -21, 47, -35, -127, -89, -109, -11, -56, 120, -118, -115, -53, -21, -8, 112, 88, 71, 110, 124, 75, 77, -92, -35, 86, -11, 47, 94, 121, 94, -39, 47, 121, 127, -45, -46, -66, 60, 51, 109, 17, 108, 88, 51, 33, 57, -114, 15, 36, -6, -38, -91, 20, -37, -95, -6, -27, -19, 15, -78, 77, 107, 112, 47, 122, 70, -11, 64, -71, -11, -72, -13, 25, 120, 118, -13, 29, -113, 21, 18, -73, -59, -34, -5, -24, 22, -110, 123, -128, -81, 81, -45, -35, 67, 0, 86, 55, -16, 0, 109, -119, 100, 62, 16, 75, -47, 84, 15, 37, -103, 81, -9, -125, 98, 39, 86, -102, -36, 122, -74, -6, 93, -112, -80, 47, -55, -28, -42, -126, 80, -63, -34, -13, -80, 51, 105, 43, 34, 20, 36, 0, 47, 123, -106, -117, -81, 118, -60, -54, -30, 34, 13, 8, 107, -62, -41, 29, -39, 48, -126, 46, -111, -3, 114, -9, -23, 125, -88, -73, 122, -48, 93, 37, 72, -32, -16, -59, 67, 63, -120, 10, -22, -81, 95, 120, -46, 102, -79, -93, 79, -43, 100, 4, 108, -112, 86, 117, 35, 36, 123, 125, 2, 116, 76, 108, -50, -82, 47, -18, -23, 92, -11, 101, 21, -93, 50, -36, 71, 32, -54, -74, -88, 76, -109, 78, 69, 41, -80, 1, 4, 61, -19, -72, -13, 111, 102, 46, 91, 93, -92, 15, 6, -120, -19, 68, -111, -45, -58, 88, -21, -30, -56, 79, 84, 44, 87, -108, 80, 88, -85, -84, 72, 87, -85, -19, -128, 100, -104, -126, -28, 85, 124, -28, -59, -10, -51, 19, 0, -100, -34, -1, -107, 28, 56, 97, -46, -43, 109, 59, 120, -114, 102, 53, -42, 42, -36, 27, -30, 79, 60, -60, 90, -8, -88, 52, -66, 62, 116, -76, -53, 75, -40, 16, 19, -21, -65, -62, 86, -38, -66, -31, -20, -72, 62, -26, 42, 110, -57, 50, -62, -110, -43, -73, 101, -44, 80, 29, 83, -94, -36, -73, -122, 112, -73, 13, -102, 115, 37, 27, -85, -96, 126, -6, 109, -67, -122, -20, -43, 102, -17, -95, -60, -120, -14, 77, -6, 120, 79, 13, -120, -121, -27, 110, -23, -92, -20, -124, -99, 20, 78, -99, -121, -51, 23, -49, 109, 91, 87, 67, 4, 82, 26, -107, 27, 65, 19, 18, 60, 50, -37, 64, 91, 35, -3, -113, 55, -93, 120, -4, 79, 105, -29, 99, 71, 64, 83, 84, 21, -35, -29, -107, 35, 95, -38, 73, 76, -105, 79, -112, 8, -116, 95, -50, 24, -55, -72, -76, 43, -8, 118, 87, 84, 95, -59, -4, -20, 115, -66, -90, -105, -95, -47, -89, 106, 66, -81, 100, -42, 68, 110, 126, -88, -1, -90, -92, 33, 72, 74, -102, 87, 102, 26, 19, -56, 121, 8, 63, -87, 127, 34, 14, 86, 112, 91, -51, -34, 24, 112, -39, -32, -50, -101, 9, 65, 73, 18, -20, -80, -85, 87, -34, 73, -3, 109, 79, 122, 92, -42, -115, 37, 26, -115, 23, -38, 68, 75, 90, 82, 108, -39, -94, -36, -62, -36, 1, 52, -38, -123, 83, -75, -59, -48, -13, 88, -56, 66, -112, 76, -14, 58, 61, -86, -15, -43, 12, 25, -111, 124, 46, 5, -47, 115, -90, 97, -101, 50, -40, -116, 86, -127, -101, 49, 48, -37, -28, -35, 13, -91, -7, -16, -42, -83, -66, -81, -36, 10, -110, -124, -77, 34, -98, 1, -55, 108, -20, 27, 67, -62, -61, -53, -87, 110, 22, -81, -56, 17, -86, 16, 34, 68, -49, 126, 51, 41, 85, 124, 116, -122, -109, -60, -79, 54, 126, 30, -16, -86, 14, -91, -83, -43, 53, -120, -13, -72, -49, -53, -11, 56, 62, 92, 43, 35, 68, -35, 114, -52, 8, -22, -3, -92, 102, -77, 36, 92, -21, 87, 49, 59, -112, 0, 20, -25, -106, 18, 46, 69, 50, -80, -71, 49, -7, -3, -47, 64, -72, -104, 121, -14, 37, -98, 95, 115, -111, -47, 82, -114, -38, 84, -29, 107, -77, 73, -20, 92, -13, -3, 123, 0, 64, 22, 0, 73, -43, -65, 103, 51, -117, -29, 28, -7, 75, 28, 90, -54, 66, -109, 102, -28, 45, 8, 31, -90, 47, -87, -2, -91, 115, -90, 67, -39, -119, 23, 113, -23, 14, 5, 56, 77, 51, 108, 93, 52, 97, 120, -63, -79, -66, 91, 124, 106, -35, 16, 28, -106, -124, -18, 35, 47, -46, -117, 109, -37, 5, -49, 4, 38, -97, 38, -57, -105, -16, -118, 105, -103, 37, -29, -40, -16, -70, -28, 53, -111, 26, -83, -116, -128, 46, 32, -49, -124, 100, 33, 48, -75, 74, 17, 24, 56, -24, -100, -61, -19, 9, 101, -22, -90, 85, -9, 2, 120, -83, 36, -82, 91, -114, 73, -40, 115, 39, -13, 34, -101, 47, 74, -51, 57, 125, 123, 85, -74, 14, -1, -62, -66, 89, 89, 79, -69, -90, -85, 80, 37, 83, 72, 48, -68, 22, -115, 1, -71, 10, -108, 38, 42, 12, -125, -122, -8, -82, 67, -51, -47, -1, -80, 90, -42, -91, 97, -63, 18, 61, 15, 125, -83, -13, -16, 8, -52, -88, 1, -57, -127, -33, 48, -47, -120, 106, 106, 120, 31, -89, -3, -52, 36, 14, -109, 52, -107, 89, 62, 105, -20, -38, -64, -77, 110, -123, -89, -22, 79, -115, -9, -37, -112, -126, -71, -87, -79, 64, -3, 43, 33, -26, 122, 114, -76, -40, 8, 11, -73, 62, -119, -95, -15, 28, 119, -38, -39, -75, 26, 57, -69, -78, -93, -43, 94, -96, -59, 83, 99, 57, 124, -8, -51, -18, 22, -113, -41, -27, -79, 16, 5, 26, 96, -114, -70, 49, 107, 84, -58, -109, -53, -104, -11, -70, 97, 65, -11, 104, 54, -34, 85, 18, 124, 47, -18, -4, -97, -124, -111, -94, 126, -103, 109, -53, -67, -102, -46, -127, -122, 79, 19, -103, 58, 120, 13, 103, -55, 19, 122, -64, 103, 27, -118, -1, -6, -5, 69, 113, -22, -124, -29, 72, 73, -45, -37, -29, -117, -80, 57, -6, -41, 74, 69, 112, -82, 31, 38, -96, -121, -119, -116, 16, -10, 93, 73, -71, -93, -23, 114, -1, -35, -103, 69, 123, 0, -122, 112, 28, 109, 120, 57, -45, 50, 98, -47, 37, 104, 7, -97, 107, 23, -74, 65, 31, 121, 78, 15, 58, -64, -103, -1, 97, -100, 123, 27, 58, -94, -103, 13, 30, -116, -17, -99, -87, 39, -44, 98, 120, -53, -65, 38, -37, 88, -107, -23, -22, 25, -31, -87, 125, 54, 91, -111, 69, 32, -95, 24, -100, 30, 92, -101, -40, -39, -93, 47, -100, -71, -22, 68, 66, -89, -36, -89, 69, -127, 58, 95, -31, 125, -31, -55, 50, -119, 74, 25, -128, 89, 21, -106, -122, 79, -61, 123, -116, -4, 64, 38, 55, -116, -76, 31, -58, 41, -40, 26, -79, 48, 59, -49, -98, -4, 95, -55, 26, -35, 11, 33, 8, 10, 110, 109, -100, -36, -95, 63, -81, 69, 108, 74, -2, 74, 67, 89, -79, -101, 30, -37, 57, -20, 101, -66, 57, -15, -42, 49, -36, -7, 76, -16, 76, -17, -15, 67, 47, 37, 115, -26, 114, -90, 83, -37, 74, -109, -100, 33, 18, -12, 119, 73, 88, -114, -107, -25, 102, -36, -27, -13, 97, -82, 115, -7, -76, -78, 121, -23, -11, -41, -35, 116, -105, -61, 93, 44, 50, 116, -95, -97, 85, 113, -118, 80, -127, -63, 117, 116, -8, 80, 23, 1, -40, 45, 70, 27, -73, 91, -110, 0, -106, 53, -110, 123, -30, -9, -33, 9, 8, 104, -57, -121, 103, -64, 14, 82, -80, -50, -25, 46, -41, -20, -14, -16, 98, -26, -123, -32, 76, 101, 16, 54, 100, -35, 114, -36, 46, -30, -82, 45, 94, -124, -30, -27, -86, -38, 83, 10, -117, 25, -44, 4, -109, 51, 104, 81, 99, -91, 64, -60, -5, 59, -43, -21, -25, -5, 33, -27, -65, -66, 110, -102, 70, -87, -110, -74, 28, -16, 74, 116, -71, -95, -61, 96, 56, 44, 85, -55, 124, 55, 63, -56, -95, -81, -83, -73, 75, 123, 71, -110, 74, -64, -76, 24, -7, -122, 112, 65, -112, -30, -74, 58, 30, 111, 76, 81, -124, 16, -30, 5, 119, -60, -3, -38, 11, 107, 72, -99, 124, 29, -28, -55, -62, -98, 87, -122, -19, -81, 95, -107, -19, 94, 125, -101, 87, 65, -110, 4, -5, -21, 69, 48, 22, 58, -9, 85, -114, -91, -29, -123, 22, 36, -45, -112, 66, 13, -50, -83, -111, -62, -58, 41, -118, -67, -84, -126, 88, -127, -42, 5, 82, -15, 71, 27, 43, -31, 106, -93, 10, -109, 12, -15, -19, -119, 33, -106, -122, 53, -78, -47, 31, 17, -105, 53, 120, -109, 80, -110, -55, -55, 79, 124, 45, 6, 66, -60, 39, -44, -27, 26, -87, -106, -55, -96, 50, 59, -58, -128, -7, 36, 90, -66, -39, -35, -94, -89, 69, -123, 66, 125, -102, -98, -63, 100, -90, -102, 61, -113, 113, -65, 109, 90, -115, -99, -83, -101, 44, 2, -83, 97, 42, -120, -54, -91, 96, -7, -17, -23, 122, -36, 15, 96, 48, 125, 40, -87, 63, -71, 110, 4, -80, 40, 25, 125, -19, 5, -23, -2, -13, -34, -123, -74, 12, -13, 27, -22, 80, 7, 122, -83, -10, -124, 62, 21, -22, -21, -104, 47, -46, 120, -55, -32, -32, -14, 119, 118, 81, 77, 78, 106, -16, -36, 37, -69, 127, -15, 46, -31, -73, -1, 34, 53, -43, 7, 33, 111, 77, 96, -102, -46, -62, -4, -83, 22, 55, -85, 122, 110, 89, 103, -7, 103, 120, -25, 46, -126, 69, -31, -4, -65, 126, -24, -5, 126, -71, 79, -94, 49, -53, -104, 99, 23, 35, 82, 8, -6, -102, -16, 74, -49, 51, -88, 9, -16, 46, -87, 43, -45, -73, 103, -111, -79, 101, 55, 80, -89, -74, -85, 121, 36, 96, 97, 50, 7, -32, 70, -87, -127, 49, 6, 41, 83, 78, 62, -54, -106, 34, -41, 59, -45, -115, -3, 35, -15, -87, 79, 83, 90, 14, -13, 71, 25, 87, -42, 19, 70, 60, 72, -93, -25, -106, -82, -96, -36, 30, -104, -36, 84, 37, 122, -125, 123, 61, -79, -99, -87, -36, -65, 105, -83, 38, 54, -84, 52, -94, -71, -100, -32, 91, 7, 8, -87, -46, 111, 59, 97, 84, 92, 88, -76, -93, -25, 25, -128, 26, 57, 21, -16, -54, -126, 35, 111, -45, 17, -9, 54, -31, 73, 42, 74, 2, 7, -13, 99, 4, -61, -32, -23, -101, -60, -21, 25, 60, 26, -58, -105, 0, 62, -8, 70, 17, -91, -52, 62, 104, 17, -16, 85, 4, -122, 16, 99, 3, -60, 108, -102, 64, -53, 123, -91, -99, -32, -98, 122, -74, 81, -36, -36, -102, 9, 82, -105, 45, -24, -104, 109, 119, 78, 124, 64, 14, -16, 90, -34, 39, -80, -24, 114, -44, -27, 29, 125, 95, -52, 34, 86, -10, 82, 53, -115, -128, 20, -124, -65, -46, 77, 62, -50, -108, -22, -77, 121, -72, 36, -65, -15, -98, 119, -92, 84, 12, 10, 10, 78, 98, -124, 31, -79, 71, 43, 10, -64, 91, 105, 61, -55, -94, 63, -46, -93, -77, -20, 27, 48, 106, -19, 99, -94, -71, 87, -96, 124, 43, -23, -126, 7, -75, -31, 67, -10, 83, -12, -62, 92, -50, 38, 72, 60, 68, 43, 93, 24, -2, 96, 7, -30, 106, 47, -40, -120, 84, -113, -23, -21, -78, -106, -89, -53, 36, 50, -13, 50, 47, 13, -36, 65, -62, 71, -54, -85, 54, -118, -128, -63, 84, 33, -49, -87, -41, -85, 50, -35, -70, 106, 76, 1, 26, 94, 54, 59, 63, -67, 92, 78, 87, 92, -16, -112, -35, 108, -94, 21, 97, -114, -51, -62, -88, 53, -64, -80, 36, 18, 31, 57, -90, 120, 20, 115, 52, 6, -44, 64, -71, -34, 49, -67, 78, -43, 99, -126, 77, -60, -2, -2, 44, 113, 83, -7, -28, 67, 102, -124, 54, 29, -105, 84, 8, 120, -11, 12, -85, 100, -43, 38, 37, 48, 15, 88, -48, 66, 98, 62, 15, 91, 109, -83, -75, -15, -16, 75, 65, -3, 43, 41, 73, 102, -94, -115, 81, -110, 127, -71, 87, 79, -40, -19, 61, -112, 64, 50, 88, 28, -47, -123, -125, -78, 79, 39, -24, -6, 59, -62, -92, -4, 114, -57, 21, 3, 39, -82, -76, -112, -8, -21, 90, -74, -52, -86, 102, -103, 123, -105, 61, 124, -62, 97, -69, -101, 50, 9, 57, 121, 23, -57, 56, -66, -69, -9, 29, -92, -12, -69, 23, 67, 16, -77, 125, -46, -44, -55, 25, -56, 108, -108, -98, 43, -64, -77, 47, -124, -123, 59, 49, 84, -70, -31, 125, 61, -14, -6, -110, 98, 57, -10, 59, 87, -77, -37, -128, 102, -22, -128, -9, 59, -18, 96, 79, -95, 87, 35, -11, 87, -45, 94, 20, 14, 117, 93, 28, -54, -28, 102, 81, 52, 98, 83, -104, 36, -109, 47, 119, -119, 101, 64, 101, 109, 72, 19, 80, 121, 22, -2, -74, 81, 121, -74, 47, -64, -73, -63, 50, -93, 40, 7, 50, 108, 124, 39, 125, -77, 21, -85, -63, -25, 47, 104, 18, 42, -124, -46, 66, 51, 112, 20, -15, -31, 70, -102, -34, -45, -62, -116, 33, -117, 42, 89, -20, -24, -79, -45, -35, -15, -90, 72, 76, -72, 99, -17, -44, 2, -115, 80, 77, -6, -24, -8, 53, 119, -111, -36, 44, 99, -86, 44, -108, 31, -18, 48, -96, 104, -55, -6, -42, -72, -112, -9, -118, 28, -37, 46, 73, 67, -79, -72, -116, 33, 75, -100, 125, 84, 114, 10, 100, 109, 52, 27, 70, 48, -82, -36, -22, -57, 127, -84, -32, 57, 118, 71, -2, 2, -112, -121, -60, 32, 40, 82, 23, -32, 44, 70, 13, 111, -85, -42, 3, 12, -7, 33, 37, 21, 58, 61, -41, -55, -105, -34, 49, 42, -75, -14, 109, 114, -93, -89, 105, 91, 58, 72, 95, 122, 13, 53, 110, -4, 36, 62, -111, -79, -79, -95, -67, -55, 125, 67, 104, 10, 9, -126, -26, -127, -105, 24, 96, -108, 85, 38, 84, 3, 65, 112, 24, -72, 67, -3, -72, -75, -66, -99, -32, 61, -49, -79, 8, -114, -15, 5, 69, 119, 55, 118, -97, 84, 126, 122, -97, 62, 22, -22, -65, -40, 0, 35, -74, -114, -127, -72, -96, -104, 41, -35, -23, -2, 95, -77, 83, 12, -7, -4, 126, -95, -57, 121, -77, 17, 26, 114, 84, 102, 91, -68, 93, -108, 103, 6, -60, -83, 111, -88, 37, -48, -108, -114, -88, -59, 40, 72, 97, 42, 116, -78, 2, 120, -32, -5, 65, 8, -108, -74, 76, -17, 117, -2, -78, 22, -37, -90, 60, -111, -106, 4, 119, 78, -40, 51, 77, 56, 89, 51, 12, 0, 117, -29, 38, -32, 73, -76, -61, -76, 106, -109, -119, -57, -104, 52, 51, -121, -36, -117, 80, 28, 71, -105, -127, 126, 23, 61, 111, -63, 4, -73, 86, -79, -81, -117, 102, -108, -91, -52, 7, -60, -38, -124, 91, 76, -3, -19, 27, -100, 2, -105, 2, -97, -7, -80, 100, 19, -35, 87, -23, -19, -79, -63, -15, -37, 22, -111, -65, -75, -98, -96, -85, 80, 13, -40, -70, 115, -109, 89, -93, 111, 8, 1, 21, 50, 108, -52, -123, -66, 5, 28, -26, -7, -11, -107, -49, 86, -103, 81, -28, 41, -24, -15, 112, -53, -91, 13, -28, 45, -80, 5, 107, -51, 31, -82, -114, 24, -123, -27, 106, 127, -27, 93, -11, -34, 47, -108, -118, -125, -19, -72, -61, 53, -31, -87, -82, 70, 122, 20, 78, 29, -1, 52, -67, 9, 25, 16, -26, -14, 94, -123, 36, 56, -70, -29, -104, -8, 24, 11, -17, 80, -79, 14, -25, 31, -118, 55, -96, -106, 1, 34, 36, 101, 115, 56, -27, -28, 2, 99, -102, -34, -86, -79, -28, 86, 17, -89, -85, 11, 8, -115, 1, -108, 80, 38, -106, -60, 114, -70, 85, 111, 47, -59, -124, -48, 103, 76, 46, 5, 95, -41, -122, -39, -72, -102, -99, 2, 70, 27, 112, 32, 7, 106, 4, 114, -107, 86, -45, -38, -8, -100, 29, 100, -128, 66, -112, -71, -47, 18, 63, 127, 4, 10, 23, -32, 107, -5, 78, -25, -53, 36, 101, 20, -68, -95, -26, 43, -21, -39, 86, -26, -119, -8, -9, -9, 90, 17, 103, 26, -84, -59, -33, 89, -27, 19, 38, 86, 27, 77, 27, -22, -22, 10, -96, -112, 77, -63, -37, 17, 123, 36, -113, 26, -122, 60, 122, 45, 91, -106, 13, -104, 84, -66, -48, -98, -10, -13, -127, 25, 0, -17, -91, 19, -80, -114, 64, -102, 29, 7, -20, -31, 47, -112, -11, -59, -97, 88, 46, -4, -52, 9, -4, -120, 75, 61, -97, -121, 63, -18, -20, 52, 45, -96, -64, 63, 45, -8, 118, 75, -107, 70, 79, 21, 72, 69, -94, 81, 63, -101, 10, 124, 20, -104, 16, -98, 58, 100, 120, 33, 44, -103, -72, -112, -53, 44, -110, 76, 1, 79, 71, 44, -22, 114, -123, -12, -110, -50, 106, -20, -111, -24, -116, 58, -60, -27, -31, -94, -10, 45, 120, 6, 71, -15, -120, -17, -89, -12, -75, -29, 119, 34, 70, 100, 57, 60, -94, -57, 95, 113, -29, -40, -94, -75, -115, -91, 17, 60, 121, -48, -37, 20, -37, -8, -90, 69, -21, -91, 84, -33, -98, -26, 98, 75, 29, -34, -37, -73, 69, 54, -18, -12, 3, 115, 76, -50, -125, 77, -8, 18, 31, 40, 15, -109, -9, -24, -126, 19, 32, 124, 56, 43, 2, -97, -92, -87, -17, 65, 70, 94, -106, -115, 19, 7, 113, -53, 37, 20, 117, 0, -75, -64, 111, -20, -78, -13, 82, 109, -105, 82, -89, 55, -101, -29, 65, -91, 44, -92, -23, 54, 31, -37, 75, -107, -41, 18, 101, 117, 120, 17, 89, 32, 58, 114, 48, 33, 74, -126, -70, -92, -30, -72, 107, 44, 119, -37, 124, 118, -36, -1, -14, -84, 96, -4, -76, -128, 117, -62, -124, -112, 12, 11, -9, 81, -78, 120, 102, -119, -56, 54, -69, 106, 10, -116, -1, 91, 32, 3, 22, 67, 101, 7, -68, -25, -24, -33, 61, 4, 64, 80, 81, -41, 63, -17, -101, -35, -59, -51, 120, -14, -61, -113, -15, -38, -10, 100, 64, 33, 46, -16, 26, -31, 22, 51, 52, -28, 53, 5, -66, 2, -41, -22, -13, 29, 109, 35, 6, -90, 71, -81, 26, -84, -111, 5, 2, 85, 125, 51, -81, -24, -39, 11, 11, -87, 101, 56, -59, 61, -119, -18, -74, 102, -124, -14, -3, -117, 8, -39, -121, 38, 36, 10, 111, -63, -101, -127, 45, -69, -105, -2, -84, 87, -126, 2, -59, 124, 66, -78, -112, 101, -48, -81, -53, -82, -52, 33, -35, -70, -95, -68, 8, -123, -87, 76, 33, -3, -105, 107, 13, 77, 117, -123, -127, -19, 11, -79, 55, -120, -120, 24, -73, 104, -25, 114, 65, -18, -18, -88, -122, 56, 91, 17, -128, 58, 43, -3, -60, 22, 20, 30, 46, 88, -73, -10, 38, 105, 45, 23, 45, -33, -37, -5, -46, -16, -1, -31, 76, 58, -52, -125, -23, 35, -35, 3, 116, 119, -43, -116, 105, -108, 53, 68, 114, -31, 91, -109, -95, 104, 89, -84, 23, -4, 57, -30, -96, 67, -48, -119, 28, 118, -120, -100, -117, 60, -73, -11, 102, -2, 120, 111, -37, -36, -110, -81, -83, 106, -75, -6, -55, 80, 35, 92, 32, 69, 16, -20, 88, 74, -43, -87, -62, 58, 118, 52, -104, 102, -121, 5, 86, 2, 104, 28, -104, 94, -63, 121, -87, 110, -118, 79, -18, 119, -15, 65, -62, -124, 4, -66, 55, -94, -51, 74, 77, 35, 14, 31, 103, 65, -19, -15, -64, -14, -62, -48, 17, -67, 58, -113, 78, 22, 94, 46, 73, -8, 23, -91, -104, 37, 69, 34, 87, -1, 115, 47, -14, -90, 121, 96, 11, -91, 84, 93, 87, -80, -112, 71, -123, -103, 13, -25, -127, 35, -122, -98, 120, 38, 86, -126, 109, 69, 79, 39, 50, -15, -126, 77, 113, -104, -117, 27, 31, -119, -88, -72, 10, 76, 0, 76, 105, -110, -56, -41, -119, -83, 106, -50, 49, -18, -48, -13, 55, 15, -39, 119, 118, -76, -29, -61, 109, -8, -31, 20, 77, -39, -67, 56, -110, -27, -28, -126, 44, -107, 39, 27, -23, -83, 23, 4, 46, 71, 90, -10, 89, 64, 77, -76, 18, -51, -15, 37, -67, -74, -39, -74, 49, 9, 92, -15, 3, -10, -94, -15, -44, 32, -50, 86, -18, -85, 55, -88, 32, -99, -79, -11, -31, 98, -11, 105, -73, 83, 10, -37, 20, -50, -51, 60, -29, 88, 81, -61, 90, -86, -2, -40, 13, 60, 116, 73, 111, 0, 25, -6, 95, 47, 111, 35, 12, -117, 98, -2, 100, 38, 123, -32, -26, 109, 64, -49, 125, -119, 94, -38, -68, 98, 91, 17, -37, 40, 107, -58, -69, -60, -36, 40, 123, -107, -92, -68, 18, -19, -35, -48, -5, 122, 10, -122, -25, 91, -114, 49, -124, 31, 27, -70, 65, -81, 112, 58, -45, 9, -30, 35, -27, -38, -20, 81, 15, 54, -12, 51, -47, -93, -20, -10, -91, 24, -27, -78, -5, -91, -81, -22, 57, 42, -40, -122, -48, 71, 75, 2, -114, 41, 109, 61, 113, 89, -97, -41, 59, 48, -107, -128, -127, 65, -5, 75, 108, 71, -85, -3, -39, -17, -29, -113, -120, 49, 38, -23, -106, 94, -118, 118, -32, 67, -104, 117, 76, -118, -26, 94, -67, -65, 65, 111, 88, 38, 112, 104, 73, 31, -9, -47, -48, 57, -37, -21, 71, -26, -60, 30, 64, 61, 109, -71, 127, 17, 35, 123, 126, -71, -91, 24, -14, 73, 28, -91, 127, 127, 26, -105, 113, -37, -90, -103, -90, 67, 0, 114, -118, 3, 87, -93, -33, 46, -39, 14, -114, -38, 31, 11, 124, -94, 59, 113, 9, 123, -57, -52, 91, -58, -84, 71, -8, 105, -46, -116, -119, 76, 38, -45, 107, -72, -120, 56, 21, -91, -38, 29, -99, 42, 16, 24, 114, 125, 22, 120, 25, -121, 39, 125, 99, -60, -2, -125, 112, -24, 23, -24, 112, 17, -104, 65, -116, 7, 5, 99, -12, -57, 102, 64, -117, -26, -48, 44, 4, 14, 32, -68, 92, 82, 81, -95, -67, 91, -116, -116, -92, -8, 40, -55, -72, -15, 80, -63, -86, 114, -115, 18, -89, -52, 108, -91, -65, 98, -29, 17, -104, 5, 85, -31, -85, 49, 52, -117, -94, 37, -45, 82, 0, -94, -106, 69, 0, -116, 7, -75, 2, 39, 74, -65, 78, -58, 69, 80, -90, -109, 49, 121, 18, -76, -65, 24, -65, 73, 13, 97, -63, -70, -82, 74, -115, -112, -65, -48, 2, -116, 121, 43, 39, 107, 91, -47, -5, 6, 66, 53, -6, 12, 98, 4, 88, -105, 103, 83, 110, -112, -88, 37, 11, -64, -98, 41, 120, -7, -49, -100, -6, -106, 64, -38, -92, -45, 62, 89, -28, -42, 14, 8, 93, 121, -1, -100, 64, -125, 39, -58, -117, 26, 36, -41, -118, -55, 100, -54, 125, -99, -22, -46, 110, 79, 26, 86, -115, 113, -61, 87, 85, 95, -30, 77, 60, -33, -16, 83, 8, 20, -114, 22, 82, 53, 57, 90, -128, 1, 55, -99, -77, 50, -54, 2, 121, -115, -122, 52, -6, 55, -96, 97, -33, -68, 63, 0, -8, -77, -23, 110, -63, 99, 23, -19, 35, -66, -105, -122, -22, -51, -115, 41, -98, 96, -16, -22, 13, 8, 97, -44, -122, 5, -5, -44, -19, -29, -83, -22, 67, -70, 59, -125, 90, 88, -53, 37, -66, -113, 94, 29, 16, -19, -115, -14, 73, -123, 123, -48, -6, -114, -21, 79, -81, 9, -112, 100, -3, -25, 57, -28, -3, 7, -11, -57, 62, -110, -44, 57, 69, -78, 48, 77, 119, -121, -3, -71, 100, 0, -108, 61, 38, 15, 90, -51, 52, -112, -62, 83, 127, 100, -84, -66, -19, 3, 119, 81, -8, 53, 34, 59, 100, 77, -22, 114, 78, -83, -23, -61, 67, -6, -101, 13, -94, 90, 76, 78, -39, 100, 32, -49, 81, -22, 15, -81, -104, 9, 53, 41, -8, -92, -124, -38, -91, -121, 43, 5, 82, -26, -15, 21, 70, 5, 126, 59, -104, 126, 63, 106, -100, 20, -77, -71, 20, -10, 100, -46, 73, -67, 80, 78, -54, 106, -12, -67, -75, 5, -70, -62, -91, -84, -22, 74, -39, 127, -117, 9, 17, -45, -7, -105, -15, 23, 32, -44, 124, 8, 94, -41, 72, -79, 96, 20, 47, 123, -50, 86, 16, -128, 49, 98, -92, 91, -39, -21, 84, -73, -85, -47, 39, 18, -14, -115, -27, 7, 92, 54, -53, -127, -54, 80, 28, -27, -54, 32, -54, -28, -100, -83, 106, 29, -30, 32, 89, -107, -52, -103, 80, -125, 124, -78, 16, 89, 26, -1, 15, 47, -121, -31, -70, -14, -22, -114, 51, 67, 117, 83, -9, -6, -110, 60, -64, 25, -60, 95, 89, 65, 89, 11, -112, -105, 127, -123, 114, -24, 52, 56, 103, -3, 7, 70, -68, 32, 107, 43, 45, 41, -27, 78, -52, 121, -17, 125, -34, -52, 37, -7, 46, -92, 47, 77, 59, 94, -76, -63, 27, 4, 109, 101, -19, -24, 39, -27, 93, -122, -119, 31, -58, -111, -44, -76, -30, 23, 25, -126, 34, -80, -35, 56, -101, 4, 120, -113, 97, 74, 43, -98, -26, -112, -65, 108, 41, 113, 124, -45, 11, -5, -77, 70, -13, -15, -14, -20, -46, 85, 120, 88, 0, 20, 70, -51, 111, -90, -25, 116, -1, 111, 100, -106, -71, 78, 117, 31, 89, -1, 0, -69, 34, 88, 3, 22, -127, -92, 112, -124, 73, -27, -7, -80, -105, 54, 82, 116, -48, 75, 76, 40, -13, 113, 35, 47, -124, -114, 107, 38, -47, 86, -95, -101, 90, -15, 90, 48, -42, 59, -120, -95, -32, 69, -105, 120, 102, 96, -63, -124, 87, 119, 8, -72, -99, 9, -90, -55, -97, 114, 107, 100, 99, -79, 59, -86, 40, 90, -81, 31, -82, -114, -78, 10, -80, 108, -87, -55, 93, 115, 80, -38, 70, -99, -110, -98, 65, -89, 105, 25, 67, -33, 29, -9, -99, 113, -57, -23, -24, -96, -121, 74, 97, -32, 11, 1, 24, 112, 123, 43, -30, 117, 15, -50, -22, -85, -13, -111, -128, 95, -49, 11, 78, -120, -16, 53, -106, 17, 91, 12, 6, 112, -95, 11, 107, -17, -32, 12, 58, 123, -124, -72, 67, -37, -85, -17, 67, -82, -109, -125, -113, 16, -75, 107, 29, 124, 84, 67, 98, -69, -12, 99, 45, 105, 120, -96, 69, 11, 42, -33, 18, 62, 65, 71, 107, 15, -67, 99, 12, 69, -66, -103, -91, 30, 75, 61, -115, -75, -63, 16, -93, -91, 1, 77, -20, 61, 20, 108, 109, -79, 62, 54, -29, -61, 80, -72, 79, 75, 36, 39, 8, 53, -83, 60, 37, -6, 3, 73, 20, -2, 28, 52, 63, -100, -120, -32, 82, -48, -14, 49, -64, 53, 73, -50, 116, -36, -123, -106, 37, 23, -27, -113, -83, 98, 86, 20, 94, -115, -82, 7, 35, 30, 64, 40, 112, 48, 95, -18, 103, -126, 7, -36, -101, 72, 107, 56, -52, 60, 106, 64, 73, -28, -106, -1, 57, 73, 104, 33, -34, 2, -42, 31, 6, 110, 33, 127, 123, 88, -32, 50, 15, 76, 61, -126, -110, 26, 39, 54, 17, -27, -55, -56, -57, 122, -35, -9, 70, -37, -72, -26, -102, -77, 7, -121, -76, 119, -111, 38, 88, 39, -1, 15, -96, -37, 127, -81, -14, -109, 120, 119, -21, -46, 121, 45, -60, -10, -28, 56, -24, 122, 15, 109, -43, -71, -91, -57, 94, -15, -127, 127, 65, 11, -119, 54, 97, -40, -72, -36, -9, -85, -80, 7, -128, 81, -119, -36, -41, -115, 77, -55, 103, -43, 6, -88, -84, 64, 1, 95, -118, 112, 106, -77, -3, -30, -22, 110, -71, -15, 65, -71, -33, -32, 127, -22, -127, 61, -53, 112, -80, 78, -91, 101, -76, 17, 60, -77, -25, -64, 50, -18, 85, 109, 79, 75, -44, -78, 97, 77, -66, 36, -7, 15, -56, -91, 92, -125, 6, 41, 45, -12, 86, 40, 25, 43, -43, -100, 68, 56, -106, -61, -73, 26, 83, 90, -5, -118, -20, -10, -13, 12, 53, 106, 105, -98, 67, 37, 32, -40, -111, 23, -42, 107, 34, -110, -69, 74, -108, 88, -5, 41, -55, -80, -62, -112, -19, 27, -100, 1, 103, 64, -84, -68, 51, 65, 118, 114, 104, 7, 80, 74, 26, 96, 19, -58, 64, -7, -85, 103, 54, 17, -79, 49, -113, -56, 112, 127, 104, -106, -122, 58, -11, -120, -41, -117, -32, -6, -104, 86, 68, -57, 46, 114, 93, 74, -119, -69, -20, 13, 103, -18, -21, 42, -85, -4, 36, -44, -93, -103, -47, -17, -18, -119, -47, 89, 117, -23, -35, -122, -114, 31, -10, 10, -34, 30, 23, -116, -105, 27, 106, 40, -109, 42, 38, -83, 98, 79, -128, -9, -27, 13, -11, 7, -50, -86, -50, 93, -27, 56, 89, -29, -16, -84, -53, 111, -109, 95, -104, 21, 62, 107, 31, 45, -82, 33, -11, -27, -25, -41, -87, 119, -110, -33, 55, 69, 22, -62, -28, 95, -91, 105, -63, -122, 111, 19, 65, -49, -73, -75, -8, 71, -22, -57, -15, -94, 44, -22, -61, 31, 7, -39, 126, -108, -63, -29, 114, -56, -91, -70, -11, -9, 42, -95, -25, -42, -116, -95, -55, 69, 77, -54, -32, -110, -33, -26, 126, 125, 108, -89, -42, 70, 36, -111, -127, 40, -84, 118, 24, 64, -21, 79, -95, 86, -14, -78, 70, -59, 61, -88, -87, -37, 113, -69, -102, -37, -56, -89, 38, 75, -27, 12, 104, -109, -55, -111, -51, -96, -102, -57, -47, 48, 32, 9, -104, 42, 59, -2, 58, 24, 39, -16, 102, -26, -72, -42, 117, -128, 62, -23, 9, -124, 30, 66, -126, -58, -70, -93, -128, -7, 60, 73, 116, -35, 56, -84, -108, -89, -22, 77, 77, -125, -100, -17, 105, -112, 58, -57, 73, -101, 74, -2, -80, -55, -41, -26, -69, 74, 80, -75, 47, 3, -94, -50, 126, -70, -30, -28, -111, -15, -42, 81, -2, 108, 44, 51, 65, 35, 121, -107, -84, 47, -72, -17, 79, 29, -42, -60, 120, 104, -34, -98, 42, 31, -62, -26, 39, -96, -127, -37, 89, 32, -58, 116, -69, -27, -11, 68, 34, 53, 25, -93, 88, 34, -54, 52, 44, -104, -70, -14, 19, 72, 118, -120, -46, 29, -125, 83, 14, 79, -3, 87, -81, -110, 104, 25, 97, -107, -31, 52, -88, 45, -122, 78, 12, 27, 99, -78, 124, -70, 121, 19, 111, 18, -31, 15, 70, 56, 126, -98, 69, 23, -83, -52, 127, -15, 50, -60, 55, 39, -113, 19, 115, -32, 98, -64, -2, 25, 14, -9, 0, -103, 60, -37, 75, -25, -52, 22, -72, -15, 12, 94, -86, -7, 107, 4, 64, 20, 86, 124, -103, 93, 66, 110, -95, -49, -116, 8, -107, 110, -10, 32, 66, 83, -48, -121, -44, 65, -66, -121, -65, -15, -99, -71, 54, -92, -25, -117, 56, -42, 94, 107, -69, -101, -57, 122, -41, 95, -18, -15, 95, -42, 10, 18, -3, -78, 84, 81, -13, -30, -18, 77, 69, 20, 21, 20, 49, 83, -5, -90, 48, -62, -85, 26, -57, 124, 86, 22, 0, 3, -23, -59, -3, -95, 48, 108, -25, -85, 18, 28, 117, 37, 125, -70, 108, -76, -100, 13, 93, 107, 43, 6, -40, 3, 98, -57, -51, 53, -128, 4, 125, -3, 57, 105, -110, 112, 123, 58, -15, -18, 73, -101, 58, 16, -54, -35, 87, -110, -80, -84, -10, 1, -116, 16, 28, -41, -120, 110, 27, -37, 58, -21, -51, -104, 64, -97, 28, -65, 77, -98, 112, -96, 108, 27, 40, 80, -53, 116, 50, -67, 25, -85, 16, 20, 60, -47, 12, -32, 88, -57, -22, -83, -59, 53, 98, 91, 67, 45, 51, -8, 19, 20, 12, 114, -12, 66, -59, -28, -38, 39, 95, 2, 126, 102, -62, -96, -101, 59, 7, -91, -53, -8, 40, 111, 96, 90, -128, -123, -25, 97, 118, 80, 86, 20, 30, -112, 14, -125, -30, -32, 122, -114, 35, 115, -73, -32, 36, 65, 101, -27, -79, 7, -122, 9, 83, -119, 54, 32, 90, 77, 11, 75, 4, 10, 25, 111, 73, -8, 127, -41, 11, 113, -24, 6, -38, -38, -106, -88, -12, 114, 114, -102, 112, -92, 65, 11, -12, 17, 86, -6, -33, 3, -57, -93, 21, 38, -4, 10, -28, -39, -16, -62, 126, 88, 29, 28, -106, -25, -47, 101, -7, 20, -60, -56, -63, 50, -73, -127, -60, 28, -113, 30, 114, -94, -2, -49, -39, 1, -28, 15, -118, 43, -98, 14, 5, -9, -113, -100, -42, 86, -80, 51, -28, 50, -47, 40, 50, -1, 77, -120, -109, 72, -91, -112, -100, 26, 30, -86, 122, -20, -96, 63, 41, 48, -100, -8, -2, 98, 90, -101, 83, 50, 84, 104, -81, -74, 24, -78, 34, 95, -12, 50, 5, -106, 47, 96, 81, 112, -117, 108, -112, -50, 28, 126, -47, -38, -90, 57, -7, -82, -112, 82, 67, 114, 118, -83, -27, -6, 122, -115, 119, -9, -2, -52, -27, 65, 9, -113, -23, -86, 10, 88, -59, 58, 47, -23, 112, -81, -57, -24, -15, -120, -83, -79, -91, -4, 96, -41, 2, 65, -95, -101, -49, -76, 111, 78, 21, -33, -62, -95, -7, 104, -54, -102, 69, -46, 17, 115, 14, -88, -37, 22, -87, 63, 48, -17, -108, 21, -109, 100, -68, -34, 116, 66, 3, 59, -97, 94, 50, 82, 127, 92, 80, -95, -54, -107, 113, 87, -26, -55, 103, -68, -3, -18, 32, 46, 63, -24, -113, -63, -81, -56, -98, 127, 65, 122, 13, -81, -121, -77, 108, -39, 45, 12, 53, -65, -14, -116, -96, 8, 14, 7, -110, 52, 125, 28, -69, 103, 35, 105, 0, 29, 109, -69, -82, 29, 30, 102, -71, 36, -76, 81, -77, -35, 7, 122, 56, -93, 60, 116, -10, -127, 17, -53, -64, -62, -108, 23, -91, -92, 91, -107, -111, 40, -72, 40, 2, -99, -78, -70, -7, -6, 18, -73, 78, 69, 57, -84, -55, -116, 59, 14, -102, 117, -110, 40, 118, -123, -50, -33, 123, 97, -93, -87, -80, -32, 110, -78, 92, -95, 123, -95, -39, -61, -12, 33, 41, 36, 9, -40, 28, 13, 28, -18, -55, 43, -50, 3, -33, -23, -20, 56, -91, -100, 0, 25, 48, -107, 113, -78, 102, 79, -6, 68, 72, 102, -33, 12, 79, -104, -6, -21, 17, 101, 123, -114, 53, 127, -128, 120, 111, -125, 1, 114, 64, 42, 119, 81, 48, -49, -128, -105, 7, -40, 96, 87, 98, -28, -18, 84, -96, -109, -94, -61, -61, 124, -99, -106, 84, 60, -59, -13, 30, -46, 81, 35, 38, -71, 71, 91, 82, -44, 74, -4, 92, 124, -9, -116, -39, 18, 24, 6, 29, -32, -117, 15, -76, 43, 23, 11, -120, 73, 1, -69, -54, 64, 18, -22, 100, 85, 49, -54, -75, -51, 120, -108, -78, 71, 90, -27, 97, -110, -24, -69, 51, -83, -102, -56, -48, -19, 91, -52, -95, -18, -112, 60, 59, -33, 126, 73, 44, -96, 114, 3, -122, 83, 32, -62, -126, -3, -27, 119, -58, -114, -99, -65, -93, 54, 109, -24, 28, 55, 60, 40, 46, -91, -56, 112, -118, 87, -50, 104, -29, -34, 123, 123, 97, 47, -108, -114, -50, -94, 70, -96, 3, -73, 126, -54, 94, 78, 40, -82, 30, 70, 91, 118, 68, -10, -78, -12, -1, -8, 75, 98, -22, -62, -123, 98, 84, 66, 122, -106, 60, 81, 92, -47, 13, -94, -34, 59, 118, -107, -63, 89, 43, 65, -55, 63, -123, -90, 108, -85, 59, -24, -19, 13, -8, -74, 104, -118, -118, 12, -74, -67, -44, -24, 94, 93, -111, -113, -98, -21, -80, 10, -89, -60, -108, -13, -27, 48, 14, 22, -31, 95, -107, -126, 107, 32, 11, 5, 20, -82, 108, 44, 94, -79, 106, -9, 73, 80, 87, 47, -27, -34, 77, -93, -94, 95, 87, -112, 39, -72, -56, 74, 19, 6, 35, -105, -15, 106, -90, -91, -3, 13, 116, -97, 69, 3, 101, 65, -39, 73, -29, -22, -24, 90, -62, 16, 116, 40, -115, -25, -4, 15, -19, -37, -32, -42, -24, 42, 45, -125, 51, -119, -74, 80, -68, 115, 91, -20, -71, 19, 75, 86, 77, -67, -12, 8, 14, -28, 87, 25, -40, 87, -14, -57, -5, -115, 27, 91, -93, -67, -67, -120, -47, -65, -78, 24, -72, 74, 74, 90, -118, 106, 103, 111, 74, 115, -27, -128, 46, 34, 80, 77, -122, 33, 124, -77, 9, -63, -75, 59, 112, 20, -37, -47, -35, -94, 63, 110, -95, 110, 27, 52, 47, 71, 3, 45, 33, 115, -46, -90, -35, 53, -7, -11, -62, 91, 43, -14, -68, -121, 30, 23, -1, 58, 106, 84, -9, -119, 59, -91, 6, -49, 2, -51, 63, 61, -22, 89, -104, 127, -92, -26, 15, -79, 24, 111, -11, 108, -112, 3, 66, -97, -103, 64, 116, 17, -35, 42, 71, 11, -84, -100, 78, 15, 89, 105, 74, 94, -40, -4, 119, -82, 37, -2, -52, -31, 45, -67, 59, -1, -117, 8, 77, 55, -91, -71, 29, -62, 2, 103, -107, -2, 99, -42, 74, 39, -96, -44, -44, -108, 92, -55, -53, -110, -120, 92, -56, 17, -44, -112, 16, 41, 75, 96, -104, -101, 97, -10, -72, 116, 15, -101, -85, 70, 43, 56, 80, 76, -29, -92, 124, 119, 8, -108, -40, -91, -84, 81, 119, 21, -43, 0, 82, -102, -60, -122, 49, -30, -70, 78, 17, -13, 100, 58, -60, 6, 92, 2, 28, -21, -115, -9, 77, -50, 75, -56, -110, 5, -126, -39, 0, 60, -115, 10, 14, 64, 93, -75, 94, -104, -71, 3, -101, -55, 15, 122, 31, 19, -63, -128, 115, -95, -9, 0, -90, 94, -15, 115, -64, -36, 23, 87, -52, -102, -111, 81, -39, -76, 3, 76, 95, -34, -3, -108, 103, -4, 37, -13, 88, 4, 37, 114, -97, -83, 66, -100, -55, -123, 37, -82, -105, -31, -102, 92, 84, 110, -35, -80, -58, -48, -2, 35, -80, 100, 80, 102, 84, -48, 7, 10, 37, -15, 5, 97, 13, 8, 75, -122, -84, 102, 51, -121, -73, 10, 84, 12, -122, 119, -116, -61, 123, 69, 95, 123, 1, 16, -24, 20, 59, 30, 102, -77, -58, -27, -63, 103, -58, 127, 10, 27, 69, -107, 44, -126, 51, -56, -74, 104, -127, 79, 63, -102, -8, 114, -62, 107, 127, 91, 18, -21, -43, -112, 125, -71, -25, -109, -6, -118, -36, -64, 4, -109, -26, -13, 28, -91, -63, -56, 41, 7, 52, 0, 35, -9, -63, 74, -56, -68, -38, -66, 43, 55, 105, 83, 105, -44, -50, -42, 41, -107, -124, 98, -114, -31, -111, -104, -9, -36, 98, -121, -16, -110, 67, 47, 74, -78, -82, 64, -121, -113, -118, -94, 69, -91, 70, 15, 27, 58, 11, -96, -115, 66, 85, -47, 48, -34, -121, -52, 31, -104, 6, 118, -3, 51, 54, -34, 108, -9, -49, -60, -7, -125, 40, -80, 40, -123, 41, 45, -101, -14, 43, 100, -68, 5, -123, 70, 125, -81, -62, 40, -47, 0, 122, 103, -27, 52, -120, 94, -95, -70, 74, 58, 0, -39, 61, 40, 88, -103, 79, 5, 6, 103, 26, -55, 27, -81, 43, 71, -86, 47, 120, 48, -121, 41, -16, -62, 12, -43, 66, 74, -98, 113, 121, 122, 63, -105, 50, -95, -6, -59, -73, 44, -75, -89, 74, -70, -80, 26, 59, 53, -37, 80, 9, -47, 108, 123, 46, 30, 49, 72, -35, -5, -67, 82, 115, 102, -46, -51, 3, -58, -61, 71, 49, 62, 93, -25, 59, 56, -29, -70, 31, 21, 83, -127, -76, -56, 28, 30, -115, 72, -30, -4, -104, 13, 67, -15, 125, 77, -24, 11, -42, -56, 95, 53, -84, -31, -15, -81, -110, 52, -72, -22, 102, -127, -80, 95, -93, -9, -120, 81, -4, -56, -123, -87, 5, 50, 108, -64, 54, 116, 98, 120, 13, -52, -5, 119, 43, -118, -17, -23, -34, 7, 100, -91, -100, -30, 64, 83, 92, -75, -55, -53, 118, -30, -75, -128, -9, -20, 66, 59, 88, 90, 119, 5, 113, 50, 5, 109, -114, -124, 27, -45, 120, 4, -41, -100, -37, -100, 37, -111, -28, 115, -111, -79, -1, -124, 84, 46, -85, 73, 1, 89, 20, -99, 18, -15, 125, 82, 56, -1, -62, -18, 59, 69, -24, -75, -87, -81, 27, -87, -59, -51, 74, -44, -118, 47, 30, 124, -105, 81, -5, -71, -72, -17, 100, -70, -39, -54, -34, -85, -14, 68, 107, -77, -38, 37, 38, 121, -73, 121, -77, -2, 52, 108, 117, -8, 31, -75, 71, -106, 47, -42, 107, -67, -126, 4, -10, -34, 55, 21, 4, -85, -120, 43, 11, -92, 43, 63, 59, -18, -56, -37, -73, -115, -1, -26, -9, 60, 31, -29, 126, 55, -70, 117, -65, 112, -86, 122, -101, -92, 64, 16, -111, 108, -32, -71, -39, -110, 44, 21, 57, -77, -47, -69, -83, -6, -49, -14, 76, -10, -56, 86, 90, -50, -20, -103, -64, 113, -28, 24, 65, 80, -39, 114, 38, 93, 31, -31, 118, -70, -64, 15, -103, -81, 87, 60, -28, -76, -90, 98, 10, -50, -2, -36, -80, 41, -26, 33, 41, 33, -122, -10, -52, 41, -91, -3, -118, -117, -91, -105, -12, 125, 87, 117, -103, 24, 119, -57, 110, -65, 124, 9, 51, -42, 78, 30, -113, -89, -123, 30, -23, -76, -36, -82, -7, 71, 36, -96, -113, -16, -95, -27, 101, 95, 88, -123, -57, 112, 37, -122, -52, 43, 120, 12, 75, 32, 110, -118, 103, 65, 34, 102, -104, -103, 8, 88, 93, 105, -97, 98, -21, -73, 120, 86, -127, 41, -58, -110, -97, 119, -92, -100, 122, 117, 16, -5, 31, -117, 47, -117, 83, 127, 15, 88, 94, -60, 2, -25, -14, -118, -116, -116, -47, 26, -6, 63, -117, -127, -68, 92, -50, -59, -23, 101, 109, -45, -32, -12, 2, 57, -84, -6, 2, -57, 76, -24, -121, -40, 18, -23, -4, -119, -53, 107, -65, 61, 91, -59, -22, 97, -36, 0, -101, -91, 68, -126, -78, -93, 55, -96, 96, -7, -86, -99, 54, 39, -96, 126, 67, 79, 15, 75, 103, 49, -48, -12, 102, 67, -104, 82, -11, 39, -107, -74, -79, 31, -19, -104, -110, -2, 0, -82, 12, -74, -63, -114, 117, -51, -102, 63, 114, 0, -39, -56, 23, -96, -63, 34, -47, -76, 76, -71, 76, 121, -90, -74, 92, 67, 18, 22, -97, 25, 38, 39, 77, 51, 76, -42, -120, -10, 94, 89, 95, -69, 57, -59, -112, 42, 60, 57, -42, -68, 119, 28, -36, 118, -124, -114, 120, -97, -81, -23, -23, 79, 110, 23, -14, -122, -25, -73, -99, 88, 70, -4, -69, -91, 118, 120, 28, -62, 49, -16, -94, -123, 126, 47, 124, 67, -70, 86, 22, -55, -42, 89, -115, -16, 104, 35, 113, 124, 88, -54, 75, 5, 61, 3, -1, 19, -86, -70, 34, 100, -49, -125, -19, 9, 100, 111, -78, -12, -41, -81, 120, 124, 127, 122, -76, -84, -47, 52, 16, 124, 2, -125, 40, 7, -22, -11, -120, 22, -68, 49, 109, 101, 116, -107, -126, -96, 96, -125, -73, -64, -3, -38, -6, -36, 20, 21, 51, 107, -102, -20, -23, 0, 31, 0, 10, -90, 103, -71, -21, 67, -59, -41, 79, 43, -51, -100, -124, 14, 14, 24, 43, 77, 123, 38, -17, -92, 38, 80, 27, 50, 18, -83, -99, -108, 97, 99, 80, 91, 85, -61, -80, 45, -114, 0, -104, 127, -40, -69, 126, -93, -2, 111, -65, 54, -82, 14, -19, -92, -96, -93, 34, -105, -57, 9, -26, 18, -28, 32, 87, -44, -76, -24, 61, -43, -88, -21, 79, -38, -5, 103, -97, 78, 99, 77, -115, 110, 100, -30, 18, 23, -101, -77, -95, -72, 119, -53, -55, -21, 90, -101, -76, -121, 23, -29, -90, -47, -10, 24, 15, 4, -40, -1, -70, -121, -65, -4, -47, 24, 11, -17, 15, -99, -45, 24, -90, 33, -36, 7, 52, 76, -104, 89, 90, -12, 6, 72, -108, -21, 97, -119, 118, -28, -123, 101, -37, 22, 127, -67, -30, 75, -47, 43, -125, 95, 25, -116, 27, -127, -53, -32, 86, 14, -121, 111, 10, -126, 71, -4, 109, 81, 98, 4, -38, -4, 70, -110, 98, 47, -99, 88, -114, -127, 99, -83, -53, 66, -34, -75, 67, 54, -71, 84, -13, -81, -8, 82, 60, -126, -38, -74, -76, 12, 31, -9, -92, 122, 122, -31, -66, -99, 114, 63, 86, 80, 72, -38, 84, -102, -40, -87, -39, -9, -108, 29, 71, -86, -20, -113, -120, 72, -57, 80, 94, -47, 89, 6, -21, 35, 65, -115, 53, 38, 40, -24, -98, 26, -37, 33, -7, 97, -7, 114, -37, -83, -47, 63, 35, 14, -112, -99, -51, 57, 122, 93, -57, -88, -4, 114, -35, 3, 79, -49, 100, -120, 88, -42, 98, 37, 106, 106, 33, -19, -111, -74, 108, 47, -57, -83, 89, 78, -2, 83, 66, 86, -66, 116, -114, -36, -60, 43, 46, 3, 5, -104, 20, -102, -50, -70, 40, -45, 32, 92, 93, -105, 120, -87, 59, -20, 85, -96, -51, 122, -81, 53, -17, -120, 16, -27, -64, 11, 35, 52, 116, 119, 122, 12, 51, 109, -26, -70, 78, 98, 99, -33, -29, -71, -14, 90, -78, -82, 77, 38, 100, 123, -109, -45, -1, -11, -82, -33, 111, 38, 21, -29, -40, 73, -45, 66, -92, 111, -48, -89, 31, -117, 79, -27, 36, -85, -49, 6, 55, 97, 54, 4, -36, 23, 68, -18, -47, -105, -34, -62, 81, 2, -14, -69, 33, 69, -43, 124, 17, 99, 107, -6, 60, 98, -92, 15, 112, 115, -73, -72, 110, 58, 99, 115, 4, 50, -39, 106, -32, 75, -55, 50, -17, -108, 102, -31, -18, 79, -43, -87, 17, 10, 16, -111, 21, -82, 19, 44, -67, 2, -111, -23, 25, 7, -19, 65, -110, 52, -60, -63, 102, 106, 27, 89, -87, 104, -38, 43, -114, 2, -49, 78, 111, -11, -13, 18, 10, 3, 120, -43, 88, 114, -110, -50, -89, -44, 76, 65, -16, -123, -106, 68, 49, -41, 107, 64, -111, -66, -4, 55, 21, 86, 2, -107, 115, 99, -89, -58, -112, 116, -127, 44, -21, 83, -128, 54, 7, 41, 12, -90, 79, -67, -89, 61, 35, 90, -21, -58, 69, 5, -13, 51, 71, 61, 25, -106, -22, -105, 86, 60, -33, 48, -9, 108, 5, 56, 41, -38, -94, -70, 22, -76, 3, 19, 42, 41, 47, 37, 80, -74, 48, 30, 127, -123, 52, -85, -5, -7, -69, -105, -99, 99, 84, 66, 42, 46, -123, 58, 69, 62, -88, 62, 122, -124, 75, -102, -85, -45, 81, 123, 33, 82, -114, 25, -90, 69, 105, -20, 120, -76, 60, 40, 10, -123, 60, -116, 26, -70, -58, -102, -65, 6, 35, -55, -103, 33, -45, -102, 33, 28, -123, 5, -18, -87, -32, -9, 28, -18, -117, 38, -20, -48, 111, 7, -111, 56, 28, 62, -1, -42, 64, -79, 67, -58, 88, 68, -75, 22, 60, -108, 104, 41, 14, 73, 105, 32, 22, -52, 35, -79, -100, 90, 33, -94, -59, -75, -37, 74, 99, -33, -38, -100, 47, -92, 66, 103, 118, -67, -95, 12, 54, 11, 91, -106, -38, 37, -18, 57, -117, -27, -102, -67, -31, 117, 76, -92, -117, 31, -122, 116, -44, -93, 45, 66, 95, -59, 92, 82, 86, -78, -19, -94, -75, 11, -77, 105, 48, -125, 78, -69, -102, -96, 15, 16, 30, -79, 84, -62, 40, 118, -96, -5, -83, 121, -92, 14, 51, 34, 96, 123, 105, -72, 36, 82, 57, -55, -58, -25, -127, 123, 34, -128, -89, -39, -71, 120, -69, -29, 18, 87, -97, 41, -76, 50, -26, 97, -98, -109, 78, -98, -54, 105, -42, 48, -78, 56, -54, -81, 119, 10, -40, 0, 63, 15, 110, -93, -66, 122, 124, 65, -9, -45, 116, 76, 80, -1, 17, 3, 113, 120, 107, -88, -94, -76, 50, 97, -6, 29, 72, 1, -1, -93, 88, -124, 99, 8, 23, 52, -3, 18, -84, -36, 48, -17, -40, -109, -9, -78, -104, 30, -124, 35, 52, -59, 41, 95, -1, 72, 96, -109, -128, -8, 69, -38, -95, 81, 121, -70, -63, -38, 80, -98, -49, -57, -54, 118, -46, -54, -19, -115, -92, -120, 55, 42, 41, -16, -76, 17, 5, -31, -83, -87, -94, -110, 95, 75, -85, 17, -75, -7, 67, -27, -2, -8, -56, 111, -103, -111, -68, -38, -53, 19, -68, 73, -66, 25, 123, 18, 64, 22, -93, -5, -18, -93, -65, 54, -15, 116, -12, 65, 24, -85, -54, -29, -9, 93, -60, -107, -14, -20, -125, -23, -11, 121, 56, 121, 25, -2, -6, -22, 5, 100, -39, 76, -27, 113, 115, 111, -18, 123, -59, 110, -98, 62, 110, 51, -6, -110, -13, 71, -40, -70, -63, 11, 91, -12, -98, -58, 64, 80, 72, -4, 100, 34, 7, 47, -9, 104, -101, 46, -92, -46, 62, -58, 9, 124, -113, -126, -72, -123, 26, -67, -47, -14, -53, 44, 100, 31, -104, -60, -97, -119, -100, -52, 60, 11, -85, -69, 7, 103, -83, -51, -112, -36, 0, -2, 36, -20, -88, -28, 26, -78, 121, -63, -114, 33, 60, 34, -55, -82, -98, 68, -108, -103, -75, -51, -55, 90, -37, 64, 13, 78, -41, 37, -73, 12, 94, 15, 94, 37, 109, -5, -65, 3, 87, 8, -90, -68, 81, 120, 75, -34, 51, 5, 82, 72, -43, -118, 23, -18, 127, 23, 4, 122, 77, 54, -2, 59, 74, -26, 18, 50, -8, 106, 107, 72, -87, 113, -103, -122, 111, 111, 47, -26, 41, -105, 99, 77, -99, -84, -71, 10, -41, -2, -86, 32, 25, -15, 58, -40, -88, -39, -6, -127, -102, -111, 2, 39, 124, 58, -88, 4, 30, -80, -119, 116, -63, 90, 109, 57, -6, -92, -88, -116, 76, -115, 125, -10, 17, -78, 119, 110, -21, 80, 120, 47, -112, 58, -122, 43, 107, -123, -107, -59, 56, -91, -6, -3, 71, -105, -66, 69, -29, -20, 51, 24, -34, 105, 61, -83, -31, 38, 26, 67, -122, 95, -103, -113, 49, -11, 80, -59, -110, 63, -89, -70, -78, -51, 34, -49, -4, 100, 104, 99, 45, 76, -111, 25, -101, -26, -80, -43, 108, 113, 121, 79, -107, -76, -123, 48, -77, 45, 30, 3, -43, 91, -42, 126, 18, 123, 80, 16, 108, 87, 126, -119, -73, -111, -40, 53, -65, -84, -31, 66, 100, -73, -4, 23, 33, 36, 89, -123, -89, -55, -62, 50, -74, -113, 17, 91, -59, 55, 30, 2, 15, -7, 26, -27, -33, 122, 77, -73, -95, -45, 115, -84, 30, -92, -90, -91, -101, -124, -83, 107, -125, 38, -5, 108, -35, 92, 73, -90, -50, 43, -74, -112, -97, -32, -84, -21, -16, -103, -37, 36, 66, -28, 0, -110, 98, -13, 11, -72, -126, -78, 95, -81, -44, -96, 90, 69, 71, -103, 8, 77, -88, 77, 36, 50, 68, -54, -16, -121, -114, -74, -95, -25, 57, -36, -67, 62, -6, 76, -39, -16, -32, 45, 95, -16, 13, -102, -8, -71, -12, -50, 34, 25, -6, -10, -114, -36, 66, -42, -116, -46, 103, 56, -14, 114, 45, 98, 89, 18, -108, 55, -67, 40, 108, 83, 105, 33, 105, -109, 31, 120, -81, 107, -119, 40, 95, 44, 56, 68, -105, 22, -80, 18, -35, 116, 93, 63, 51, 124, 96, 82, 123, 62, 125, 108, -33, 51, 77, -36, 57, -119, 52, 70, 64, 43, -64, -44, -108, 65, 73, -13, -125, 105, 127, -88, -41, 103, 79, -43, 15, 109, 125, -89, -127, -121, -87, -38, -41, 32, 32, -94, 91, 74, 95, 41, -20, -35, -61, 74, 75, 27, 70, 45, -20, -96, 17, 69, 52, -108, 8, -37, 119, -53, 41, -111, 108, -52, 16, -54, -34, 49, 17, -100, -107, 72, -110, -73, 84, -89, -47, -108, 20, -12, -42, 126, 37, -19, 60, -79, 36, 34, -70, -100, -64, 99, -83, 31, 2, 119, -21, 118, -127, 77, -102, 3, -17, -61, 95, 80, -96, -87, 61, 59, 90, -88, -105, 77, 12, 16, 24, -71, -114, -10, 22, -28, 124, 99, 120, -68, -91, -111, 114, 67, -27, 94, 2, -24, -84, -120, -23, -107, -38, 3, -52, 65, -14, -67, 28, -103, -126, -72, -15, -111, -68, 86, -106, -92, 40, 70, -40, -31, 96, -58, 0, 58, -66, -71, -28, -124, -5, -92, 19, 89, -102, 101, -119, 94, -88, 87, -62, 108, 106, -64, -108, -127, 76, -119, 80, 101, 119, 52, 76, -93, -128, -108, -13, 35, -20, -48, 41, -91, 81, -4, 116, -90, 121, -100, -100, -77, 23, 90, 56, -41, 111, 103, -48, 125, -24, 51, 110, 107, 96, 47, 79, 24, 67, -9, 68, -91, 82, 67, -100, 92, -17, 52, -16, -5, -2, 40, 26, -46, 108, 72, -86, -88, 82, -52, -84, 21, 4, 77, 59, -70, 27, -60, 84, -10, 43, -10, -51, 29, -14, -37, -99, 70, -32, 1, 52, -46, 122, 112, 51, 19, -67, -100, -78, 24, 118, -81, 5, 93, -114, 46, -47, -76, -86, 127, -34, 107, -49, -57, -114, 96, 119, 75, 45, 93, -61, 53, 2, 78, -9, -59, -38, 11, -52, 126, -118, -39, -111, 39, -52, 75, -25, -45, -116, -20, 93, -128, 23, -48, 0, 127, -118, 10, -34, 113, 25, -84, -40, -114, 88, 33, 34, -28, 102, 120, 73, 109, 18, -123, -53, -30, 11, 72, -68, -123, -66, -17, -26, 113, 38, -107, -101, 114, -12, -106, 127, 19, -22, -128, -27, -29, 92, 62, -76, 45, 97, 69, 48, 12, -8, -80, 71, 67, -78, -118, -91, -102, 88, 15, 100, -128, -23, -126, -77, 71, 62, 107, 11, -67, -84, -106, -75, 58, -25, -35, 55, 33, -65, -128, -42, 22, -102, -14, 26, 71, -30, 108, -1, 72, -36, -93, -45, -124, 43, 122, -105, -81, 4, 1, 102, -55, 68, -113, -24, -33, 34, -82, 123, -10, 48, 103, 78, 70, 50, 77, 34, 86, 62, 33, 37, 81, 76, 53, 20, -83, 75, 45, -60, 68, 72, 65, 93, 89, -6, -112, 43, 82, 94, 2, -22, -104, 12, 55, 50, 13, -39, -95, -70, 71, 23, 31, 39, -35, -9, 83, 9, 99, 14, 1, -38, -84, -115, -58, -3, 90, 6, -68, -124, 123, 90, 43, -80, -84, -84, 103, 32, 44, 70, 58, 56, 75, 117, -116, 106, 111, -119, 101, 89, 27, 109, -92, -17, -53, 47, -37, -43, 3, -50, 59, -43, 115, -128, 110, -80, -40, 113, 38, 107, -82, 17, 12, 2, 47, -8, -12, -24, -54, 112, -16, 78, -90, -109, -82, 60, 115, -43, 127, 33, -109, -88, -28, 102, 92, 91, 16, -53, -31, 89, -63, -45, 22, 27, -25, -69, -113, -116, 25, -112, 37, 69, 110, -66, 93, 60, 25, -66, 6, 57, -48, -10, -87, -51, 10, -65, 124, 100, 25, 58, -45, 64, 127, -113, -126, 59, 44, -95, -122, 91, 99, 92, -78, 3, -96, -93, -102, -73, 23, -42, 60, 89, 31, 112, -18, -83, 6, 125, 29, -83, 54, 111, -2, -83, -124, 25, -56, -102, -67, -20, -40, -64, -120, 9, -84, -64, 127, -4, -21, 54, -98, -42, -96, -126, -65, 78, -33, -88, -81, -62, -63, 58, 24, 66, -24, -94, -74, -15, -107, 72, 14, 66, 18, 17, 56, 35, 45, 96, 29, 20, -127, 40, -44, 48, 82, -51, -14, -108, -71, 126, 2, -38, 82, 28, 6, -27, 57, -39, 109, -30, 49, -84, 35, 87, 38, 106, -90, -99, 115, -67, 100, 0, 1, -66, 71, 63, -28, -57, 28, 6, -105, 88, 8, -61, 5, -27, -53, -112, 85, 68, 86, 122, 4, -81, -63, -50, -45, -74, 90, -78, -24, 46, 10, 72, 14, 29, 64, -101, -128, -73, 90, -16, -14, 13, 124, 12, 59, -96, -32, -10, -35, 116, 90, 61, -101, -56, 73, -96, 71, -41, -49, -39, 68, -126, -124, 59, -82, -73, 102, -12, -114, -14, 63, -15, -89, 121, 46, -112, 15, 78, -43, -60, 36, -67, 22, 106, -10, -49, 1, -14, 49, 46, -16, 35, -81, -4, -49, 41, 45, -92, -34, -54, -118, 52, -42, -9, 99, -14, -108, 57, 73, -14, 112, 122, 66, -128, 27, -90, 80, -26, -74, 30, 90, 48, 25, 64, -66, 75, 74, -85, 50, 60, 47, 106, 88, -124, 47, 101, -109, 4, 18, -11, 72, 91, -105, 112, -14, 121, 127, 75, -96, -65, -58, -11, -64, -40, 51, 93, -114, -1, 23, 18, -78, 46, -46, -37, 50, 28, -107, 57, 122, -54, 9, 7, 76, 11, 122, 58, -17, -114, 125, -10, 54, 8, 46, 84, -125, -124, -5, -56, -29, 11, -108, 14, 94, 103, -49, -39, 73, 74, -70, -83, -13, -12, 18, -89, 109, 97, -100, -34, 86, -80, 5, 12, 124, -64, 93, -72, 36, 123, 69, 41, -58, 82, -114, 43, 96, -123, -121, 21, 25, -100, 99, -53, 90, 119, -87, 15, 95, -84, -98, 11, -15, 108, -111, -15, 76, 84, 123, -116, 63, -24, 2, -121, -33, 78, 92, -109, 116, -65, -15, 9, 49, 85, -17, -28, -48, 97, -48, 70, -102, 8, -49, -101, -115, -32, 88, 80, -105, -4, 123, 26, -29, -54, -102, 89, 50, -13, 105, 84, -65, 53, 113, -106, -59, 9, -86, 95, 26, 74, -121, -70, 32, 45, 22, -106, -128, 80, -57, 41, -123, -11, -23, -125, -70, 50, -104, -12, -109, 30, -5, -20, -52, 62, -68, -88, 13, -98, -9, 6, 94, 97, 36, 110, -52, -19, 83, -7, -54, -45, 45, -23, -90, -98, -98, 79, 84, -67, 85, 2, -10, -78, 24, 56, -29, -40, -33, -40, -26, 48, 7, 101, -45, -41, 115, 24, -26, -63, 29, -58, 52, 58, 69, -36, -80, 75, -21, -93, -110, 89, -77, 48, -122, -25, -115, 7, -96, 91, -71, -23, -16, -59, 22, 121, -74, -89, -97, 49, -77, 33, -63, 39, 3, 59, 109, -59, 109, -94, 123, 4, -110, -127, -38, -11, 92, -18, 66, 67, 58, 56, 53, -107, 16, 107, -78, 52, -73, -94, 6, 34, -85, 76, -112, -94, -90, 58, -40, 37, -3, -77, -90, -102, -1, -79, 4, 38, 27, 111, -109, 8, 18, 120, -80, 3, 99, 5, -128, -62, 97, -27, 110, -111, 23, 74, 80, -92, -108, -17, -115, -83, 59, -3, -122, 37, -118, 54, -18, -88, 120, 67, -25, -87, 77, -35, -34, -14, -43, -58, 99, 115, 40, -85, -100, 79, 63, 115, 75, -48, 55, -20, 41, -75, -50, -27, -93, -2, -9, 35, 35, 75, -39, 109, -60, -73, -10, -62, -128, 90, -66, 13, -79, 74, -14, 108, -36, -89, -46, -45, 111, 0, -68, -14, -106, -5, -12, 52, 35, 10, 0, -1, 77, -14, -59, -54, -29, 34, 123, 116, 99, -32, -109, 15, -125, -78, 35, -119, -89, 81, 59, -116, -110, -70, 96, -22, -16, -38, 97, -35, 56, -61, -126, -103, -13, 85, 96, -7, 68, -113, -77, -105, -30, 0, -45, 69, 68, 32, 22, -117, 43, -46, 18, -94, 114, 37, 35, 94, 125, -52, -16, 15, 118, 25, -108, 118, -49, -126, -125, 27, -83, 95, 62, 2, -63, 95, 94, -54, -9, 82, 51, 28, -29, 46, 60, -4, 90, -86, -118, -74, 91, -63, 127, -104, -32, -2, 120, -69, -22, 28, 7, 101, -42, 95, 99, -127, 113, -89, -119, -89, 81, 50, -53, -3, 118, -35, 2, -23, 18, -19, -99, -96, 102, -114, 26, 75, -113, -4, 53, 95, -36, 18, -4, -64, -112, 49, 75, -73, -102, -58, 5, 64, -43, -25, -37, -1, -110, 44, 92, -85, -124, -128, 30, 3, 24, 71, 26, 107, -112, -37, 53, -113, 126, -35, 19, -53, -46, 83, -37, 70, 78, -109, -15, -85, -30, 3, 92, -92, -65, -109, -35, -96, 32, 105, 126, -13, 126, -89, -16, 74, -113, 23, -128, 85, 45, -11, -36, 9, -1, -38, 106, -109, -33, 80, -94, 85, 127, 56, -72, 116, -119, 76, 63, -123, -13, -103, 65, -2, -70, -70, 40, 87, 40, -103, 96, 23, -43, -69, -74, -30, -56, 125, 72, -42, 11, 71, -32, -6, 95, -40, -14, -12, -71, 119, 26, 13, 32, -80, -126, -58, -76, 107, -6, 15, 110, 13, 107, -36, -118, 36, 0, 89, 108, 53, 63, -68, -80, -38, 61, 59, -120, -6, 42, 39, 114, -38, 26, 85, 125, -120, -113, 101, -30, -43, -29, -65, -85, -41, 12, 9, -38, 100, -26, -29, -30, 95, -66, 88, 56, -61, -79, -78, -119, 124, -92, -10, 22, 67, 103, -27, 98, 9, 13, 87, -122, 59, 114, 6, -55, 59, 30, -5, 53, -76, -117, -86, -14, -13, -45, -92, 40, -16, -9, 52, 71, -65, 56, 97, -78, -100, 16, 39, -24, 117, -62, -126, -39, 108, 49, -88, -112, -13, -63, 56, 111, -45, -124, 96, 31, 14, -105, 23, -117, 11, 65, 23, 99, 27, -51, 73, 126, -44, 82, 23, -47, 17, -86, 92, 27, -27, -87, 47, -99, 21, 45, -8, -127, 88, 56, 102, 9, 83, -52, -104, -30, -9, 48, 116, -17, -69, -53, 75, -20, 86, 1, 80, -89, 56, 17, -81, -62, -99, 11, -7, 99, 108, -32, -21, -27, 92, 79, -98, 44, -61, -3, -106, 31, 57, 104, 88, -91, 36, -11, 79, 89, 126, -27, -124, 25, 9, -69, 125, -105, -29, 38, -99, -30, -60, 36, -52, 15, -104, 58, -122, -68, -101, 85, 25, 45, -128, 21, 30, 19, -81, -99, 34, -87, -79, -23, 58, 21, -108, 33, -124, -47, -46, 88, 96, -90, -28, 49, -116, 19, -56, -72, -43, -95, -120, -13, 6, -100, 26, 11, -72, 51, -100, -104, 64, 75, -21, -6, -127, -113, 9, -2, -92, -61, -24, -118, -91, -27, -53, -105, -69, 127, 109, 85, -126, 126, -66, -98, -83, 45, -44, 117, -120, 17, 108, -117, -7, -71, -78, 70, 48, -47, 74, 55, 69, -15, 0, 54, -92, 99, -109, 7, -9, 48, 106, -75, -26, 27, 26, 70, -63, -26, -75, 44, -81, -44, 0, -111, 83, 12, -116, 9, 58, -58, -14, -74, 8, -33, 0, 107, 65, 22, 84, -49, 36, -36, -12, -53, -40, -5, -114, 97, 84, 81, -2, 41, -41, -69, -110, 125, 31, -8, 57, -3, -96, 124, -12, -91, 7, -33, 15, -82, 20, 47, 10, -96, 67, 3, 3, -44, 77, 78, 63, -101, 2, 81, -5, 79, 21, -34, 79, -30, 106, 68, -95, 5, 120, 36, 24, 81, 5, 41, 74, -31, 117, -7, -23, -47, 114, 80, -8, -35, -122, 100, -8, -45, -79, 8, 96, 4, 105, -16, -94, 79, -36, 4, -53, 61, -99, -112, -69, 117, 69, 99, -7, 10, 13, 98, 60, 10, -2, 112, -112, -43, -79, 82, 47, 117, -116, 100, 77, 122, -57, -124, -63, 33, 42, 126, 58, -86, 97, -68, 61, -95, -79, -53, -27, -26, 48, 92, -42, 4, 98, -18, -110, -91, -64, -64, -10, -121, -50, -40, 104, 13, 75, -60, -107, -47, 95, -57, -58, -97, 66, 62, 116, -91, 125, -24, -112, -103, -17, 35, 80, -81);
    signal scenario_output : scenario_type := (-54, -36, 49, 127, -29, -76, 13, -12, 96, -59, 3, 18, -52, 10, -74, 106, 112, -58, -107, 54, 64, -116, -66, 36, 65, -3, -13, -44, 69, 127, -117, -39, 88, -18, -111, 79, 69, -38, 65, -123, -81, 52, -37, 80, 64, -63, 17, 54, -33, -73, 38, -36, 18, 86, -128, 37, 109, 16, -59, 3, 90, -88, 21, 53, -103, -111, -18, 112, -33, -13, 87, -52, -43, 59, -10, -90, -10, 124, -16, -122, 127, 8, -112, -36, 127, 7, -128, 29, 116, 81, -122, -50, 121, 63, -93, 16, 45, -3, -93, -22, 13, -45, 119, -68, -64, 3, -7, 2, 78, 106, -128, -52, 7, -18, 85, 59, 21, -96, -108, 93, 39, 43, 22, -98, -48, 60, 98, 8, -69, -12, 3, 57, -39, -122, 0, 43, 114, -36, -55, 11, -32, 16, 3, 21, 95, -97, 8, -10, -22, 127, -60, -11, -57, 50, 17, -87, 100, -13, -5, -2, -6, 36, -101, -44, 0, -11, 48, 44, -10, -70, 11, 70, 86, -95, -128, 127, 88, -128, -80, 43, 18, 24, -18, 49, 1, -22, 48, -66, 22, -28, 78, 55, -107, 68, 71, -23, -31, 24, -28, -63, -1, 47, -70, -31, 5, -36, 81, -29, -47, 55, -5, -11, 76, 57, -87, -85, 118, 3, 12, 54, -128, -73, 127, 16, -128, 96, 96, -22, 49, -118, -38, 127, -81, -98, 69, 107, 10, -112, -106, 93, 108, -100, -1, 44, 7, -5, 6, 36, 6, -16, -95, 59, 64, -57, -39, 27, 98, -38, -128, 0, 114, 15, -44, -95, 34, 27, -7, 127, -128, -60, 127, -38, -48, 80, -106, -49, 0, 78, 12, -23, 124, -128, 1, 28, -108, 57, 38, 2, 18, 13, 48, 39, -64, -128, -8, 108, -66, 31, 44, -39, 95, -13, -50, -13, -42, 12, -38, 13, 127, -24, -128, -50, 3, 32, 21, -47, -32, 127, 76, -113, -60, 66, 127, 5, -128, 33, 59, -128, 0, 106, -54, 33, 102, -50, -128, 7, 127, 50, -55, -118, -31, 27, 33, -50, -31, 112, 12, -33, -13, 3, 28, 0, -63, -63, 36, 102, -5, 2, -24, 0, 36, 37, -45, -117, 57, 27, 16, 24, -11, 24, -36, -118, -31, 127, 15, -39, 28, -48, 75, -7, -7, 43, -71, 5, 38, 2, 43, -63, -48, 37, -10, -23, 27, -64, -93, 52, 69, 54, 55, -29, -29, 57, -78, 6, 11, -69, -34, 75, 80, -36, 21, 38, -100, -69, 113, -76, -100, 31, 71, 63, 39, 28, -128, -21, 95, -54, 43, -47, -24, 111, -100, 42, 95, -29, -32, 22, -42, -58, 7, -59, 13, 117, 43, -127, 79, -32, -113, 127, -29, -58, 80, 5, 44, -32, -128, -13, 127, 6, -128, 50, -13, 42, 127, -128, -124, 117, 27, -69, 11, -7, 43, -34, 1, 32, -15, -28, -11, 3, 17, 93, 38, -75, -92, 127, -36, 3, 15, 0, 50, -107, -50, -7, 121, 53, -118, 52, 127, -69, -102, -57, -34, 127, 58, -18, 16, -80, -11, 29, -32, 8, 17, 39, 27, 12, 10, -128, -13, 31, 86, -26, -60, 0, -43, 58, -38, 111, -16, -36, 31, -48, -2, -85, 79, 100, -43, 16, 8, -58, -75, 43, 127, -64, -87, 103, 86, -128, -128, 39, 109, 32, 0, -16, 15, -45, -128, 33, 64, 49, -55, -3, 73, 22, 24, -113, -101, 69, 121, -45, -128, 98, 127, -91, -92, -17, 50, 88, 13, -98, -68, 49, 32, 28, -38, -54, -10, 50, 0, -42, -5, 12, -10, -24, 3, 0, 2, 97, 18, 15, 64, -128, -43, 112, 38, 27, -127, -21, 127, 29, -55, -43, -64, -90, 71, 7, -69, 24, 88, -8, 11, 31, -68, 28, 101, -36, -66, -3, 16, -3, -8, 3, 34, -26, -117, 47, 47, -21, 74, -45, -32, 88, -57, -50, 69, 2, -96, 117, -27, -59, 127, 5, -31, -71, -53, 114, 86, -85, -74, -52, -22, 101, 17, -15, -16, 31, 23, -37, 81, -52, -79, 37, 32, 11, -11, -5, -80, 75, 2, -128, 74, 107, -32, 24, -17, -57, 42, -27, -39, 39, 37, 15, 55, -108, -87, 53, 12, 54, 74, -64, -117, 21, 107, -38, 15, 24, -128, 88, 75, -128, 38, -11, -58, 64, 11, -65, 42, 3, -59, 6, -13, 119, 65, -3, -71, -47, 127, -28, -112, 44, -29, -34, 29, 23, 16, 54, 2, -8, 8, -97, 7, 42, -79, 74, 95, -68, 28, -6, -68, 22, 28, -15, -58, 11, -5, -81, 34, 68, 16, -23, 15, -27, -37, 109, -6, 0, 91, -23, -96, 11, -21, 34, 63, -58, 0, 39, 2, 1, -32, -66, 68, 0, 16, 50, -24, -52, -103, 55, 113, 16, -108, -128, 44, 69, 97, -78, -18, 127, -128, -109, 98, 102, -66, 0, 124, -128, -96, 50, 47, 2, -86, -29, 27, -24, 18, 91, -45, -34, 0, -34, 24, 47, 54, -93, 15, 29, -75, -12, 100, 101, -63, 48, -80, -85, 127, -78, -73, 85, 26, -7, -80, 80, 13, -34, -21, -114, 127, 65, -87, 11, 87, 16, -114, -15, -22, -10, 6, 0, 65, -8, 75, 49, -43, -118, -7, 102, -86, -27, 127, -7, -78, 44, -6, 54, -44, 1, -24, -16, 63, -71, 64, -52, -96, 127, 122, -65, -100, -22, 3, 3, -44, 34, 60, -22, 79, -8, -17, 48, 21, -57, -48, 54, 16, -87, 27, 101, -58, -87, -3, 49, 3, 15, 16, 57, -113, -49, 75, -59, 0, 13, 7, -33, 37, 16, -102, 5, 127, -60, -22, 127, 2, -17, -18, -21, -103, 68, 33, -128, 17, 111, 32, -63, 24, -33, 42, 24, -65, -22, -23, 60, 23, -38, -39, -21, 57, 42, -92, 80, 65, -103, 28, 2, -57, -34, 42, 10, 7, 76, -122, 0, 75, -53, -55, 98, 45, -11, 81, -122, -74, 10, 65, 12, -66, 26, 29, -22, 39, -44, -107, 113, 50, -63, -70, 111, -5, -128, 90, 88, -71, 10, 15, 26, -16, -45, 33, -24, 44, -39, 3, 93, -87, 18, 90, -128, 2, -11, 36, 116, -111, 11, -24, -76, 121, -44, -26, 78, -13, -24, 57, -17, -26, 60, -27, -96, -17, 111, -59, -7, 109, -48, -52, 86, 66, -44, -11, -88, -86, 50, 109, 85, -128, -49, 93, -85, 81, -29, -15, 127, -71, -57, 69, 13, -114, -64, 71, 31, -8, 50, -29, -2, 2, -1, -44, 32, 5, -39, -29, 24, 127, -45, -128, 47, 127, 21, -57, -63, -28, -24, 87, 10, -60, -66, 44, -6, -18, 127, -37, -101, 113, -22, -17, 108, -3, -111, -79, 45, -18, 6, 48, 79, -49, -96, 98, 63, -128, -63, 5, 54, 114, -6, 23, -27, 18, -48, -57, -2, -92, 58, 102, -11, -65, 93, -17, -22, -34, 33, 80, -42, -87, 42, 127, -124, -60, 15, -32, -47, 80, 42, -21, 50, -96, 65, 45, -70, 2, -64, 31, -6, 57, 2, -70, 17, -33, 32, 10, 90, -13, -87, 26, -8, 31, 86, -21, -22, 5, -93, 0, -26, 50, 37, -65, -8, 44, -42, 65, 74, -28, 16, -88, -65, 108, -7, -31, 37, -2, 3, -90, 10, -8, 79, -15, -42, 18, 8, 54, 31, -1, -128, 45, 123, -54, -22, -8, -57, -53, -5, 28, 15, 88, 96, -100, -128, 127, 44, -121, 55, 107, -103, -52, 93, -63, -12, 68, 23, 8, -5, 33, -74, -29, 53, 37, -26, -128, 47, 22, 42, 92, -43, -128, 87, 8, -128, 45, 27, -31, 90, -13, -10, 121, -13, -103, -112, 127, 58, -128, -28, 127, 31, -71, -57, 76, -50, -1, 116, 1, -66, -11, 109, -128, 0, 127, -54, -128, -65, 71, 13, -73, 68, 71, 63, -87, -38, 95, 15, -123, 33, 52, -112, 29, -32, -24, 70, 65, -75, 53, -8, -48, 127, -39, -85, 96, -27, -128, 112, 18, -1, -12, -128, 100, 33, 22, -45, -38, 49, -17, -8, -2, 108, 22, -8, -44, -16, -87, 31, 127, -53, -52, -10, -74, -54, 34, -12, -34, 22, 12, 96, 73, -123, -3, 34, -65, -38, -6, 101, 29, -101, -52, 101, 97, 7, -59, -63, -24, 26, 2, -50, 37, 31, -18, 93, 27, -102, 18, 38, 53, -38, -38, 80, -23, -42, 16, -32, 47, -29, -113, -11, 42, -8, -24, 88, -11, 31, 43, -5, 8, -52, -70, -59, 87, 37, 55, 6, -93, 65, 45, -26, -29, 0, -23, 66, -73, 2, 127, -128, -15, 88, -79, -11, -3, -42, 66, 36, -96, 87, 10, -127, 70, -18, 42, -5, -43, 26, 75, -29, -74, 127, -73, -100, 8, 80, 87, -128, 32, 95, -128, 68, 117, -116, -8, 50, -22, 74, -81, -38, 85, -44, 38, -29, -116, 13, 43, 8, -3, 12, 0, -92, 91, 127, -15, -128, -7, 117, -26, -50, -22, 27, -68, 39, 98, -70, 6, -17, 57, -3, -12, 50, -128, 10, 100, -103, 36, 127, -128, -1, 27, -58, 13, 34, 49, 16, -45, -88, 127, 26, -74, 75, -66, -128, 107, -1, 3, 127, -116, -16, -5, -27, -10, 74, 23, -128, 44, 54, -55, -59, 86, 1, -49, 0, 65, 122, -73, -38, 58, -75, 1, -1, -34, 127, -29, -32, -2, -52, 78, 55, 24, -102, 26, 10, -119, 26, 91, 18, -52, -33, 7, 86, 0, -109, -65, 50, 5, -45, 117, 43, -80, 95, 18, -128, 65, 70, -32, -78, -22, 76, 21, -60, -86, 33, -16, 98, 7, -128, 111, 112, -102, -112, 108, 52, 28, -78, -23, 127, -49, -119, -91, 70, 112, -24, -1, -12, -39, 78, 18, -73, 57, -10, -98, -38, 59, 96, -103, -52, -11, 113, 10, -122, 107, -3, -5, 10, 0, -24, -65, 101, -26, -45, 127, -50, -7, 8, -128, 91, 112, -112, 0, 44, -45, 21, 48, 31, -100, -15, 101, -12, -32, 36, -52, -24, 27, -98, 70, 29, -13, 106, -22, -10, -88, -7, 21, -48, -5, 70, 69, -29, 71, -123, -24, 65, 17, -57, -90, 58, 60, 88, -128, -42, 12, 18, 127, -42, -36, -70, -22, 127, 8, 15, -15, -124, 13, -18, -59, 59, 111, 78, -52, -128, 0, 127, -21, 13, 59, -86, -113, 75, 124, -34, -90, 16, -44, -86, 23, 6, 52, -13, -27, 124, -1, -113, 13, 32, -27, -24, 66, -6, -85, 21, 45, 93, -47, -2, -32, -54, 42, -81, 78, 2, -68, 31, -7, -16, 31, 68, 16, 47, -29, -128, 60, 16, -91, 127, -16, 0, 44, 3, -50, -39, 50, -8, 59, 13, -70, -28, -34, -57, 29, -18, 86, 55, -23, -76, 22, 127, 7, 3, -36, 12, -87, -103, 127, -33, -24, 34, -97, -39, 123, 66, -15, 69, -73, -93, -27, 118, -5, -128, 49, 42, 54, -68, -37, 34, 60, -38, -81, 88, -33, -58, -7, 97, 74, -47, -95, 39, 88, -8, 48, -29, -98, -31, 27, 48, 50, 47, -111, -18, 15, -17, -12, -48, 0, -18, 91, 127, -55, -98, 111, -3, -45, -12, -68, -3, 0, -21, 64, 122, -15, -18, 6, -32, -54, 17, 121, -90, -32, 98, -24, -15, -88, 36, 5, 34, -2, -64, 24, -60, 93, 39, -31, -7, -50, 93, -60, -103, 81, 58, -81, 34, 6, 1, 33, -55, 123, -97, 1, 127, -118, -90, 60, 42, -3, -29, 37, 13, -52, 23, 37, 8, 0, -11, -63, 44, 85, -17, -102, 23, 22, -21, -63, -18, 63, -70, 53, 76, -17, 29, -100, -73, 127, 43, -71, 27, 7, -73, -29, 63, -34, -66, 65, -22, -48, -32, 127, 127, -55, -3, -54, -127, 18, 80, 66, -28, -1, 66, -27, -91, 54, 39, -38, 28, -11, -12, -60, -34, -17, 10, 36, -26, 50, -36, 5, 69, -28, 3, 52, -71, -6, 57, -121, 49, 3, -48, 10, 98, 34, -93, 15, 85, -24, -92, -18, -10, 88, 76, -90, -34, 34, 26, -48, 7, 123, -128, -49, 54, 52, -26, -128, 127, 106, -128, 49, 90, -128, 11, -16, 29, 22, -37, -6, -10, 73, -96, 3, 39, -23, 47, -42, 21, 98, -97, -80, 127, 45, -100, 1, -24, -16, -12, 52, 3, 36, -21, -53, 45, -28, 3, 64, -16, -3, 31, 7, -75, 3, 34, -52, 127, -36, -128, 39, 63, -22, -17, -43, 10, -16, -28, 38, -1, -55, 93, 117, 0, -96, -109, -6, 97, 50, -57, 71, 96, -55, -91, -34, 44, 113, -108, -47, 73, 0, 6, -64, 71, -3, -36, 100, -38, 21, -78, -5, 50, -59, 55, -16, 18, 13, -88, 60, 12, -31, 91, 29, -96, -98, 60, 107, -97, -95, 37, 68, -16, -60, 43, -32, 21, 95, 16, -49, -28, -74, 13, 127, -78, -49, 70, -97, 58, 47, -2, -37, 23, 13, -45, -13, -57, 90, -12, 57, -1, -121, 75, 16, -111, -31, 13, 119, 34, -58, 49, 48, -91, -90, 5, 88, 96, 10, -102, -65, 10, -24, 12, 87, 1, 26, 12, -28, -5, 26, -7, -97, 13, 96, 81, -85, -8, -43, -22, 80, -44, 32, -58, -31, 127, -103, -12, 64, -88, 16, -49, 57, 88, -52, -10, 16, 64, -38, -26, 88, -11, -113, 8, 121, -95, -128, 2, 32, 127, 7, -23, -16, -50, 103, -34, 3, -8, -107, -2, 43, 81, 12, 34, -121, 27, 127, -68, -109, 66, 55, -65, 65, 52, -29, -22, 18, -93, -37, 22, -29, 54, -52, -100, 127, 91, -63, -32, 59, -43, 21, 108, -70, -59, -81, 39, 95, 15, -33, -88, 60, 78, 6, -8, -123, 36, 111, -117, -91, 31, -23, 29, 108, -1, -55, 63, 38, -64, 34, -23, -49, 6, -69, 86, 111, -106, -100, -21, 95, 113, -17, 0, -23, -8, -55, -88, 85, -28, -49, 98, -26, -27, -17, -26, 91, 13, 36, 70, 1, -1, -128, 23, 13, -48, 116, 17, -18, 11, 64, -128, -90, 127, -21, -128, 45, 1, 34, 63, -128, 66, 12, -78, 127, 8, -74, 16, -38, -76, 49, 127, 0, -121, -59, 75, 63, -24, 48, 39, -112, -42, 75, -50, -60, -27, 95, 49, -95, 79, 92, 1, 5, -78, -50, -33, -59, 100, 98, -27, -128, -8, 91, 63, -57, -128, 43, 127, -79, -90, 21, -64, 27, 102, 2, -101, 69, 43, -107, 13, 127, -71, -86, 127, -32, -59, -23, -33, 70, -1, 36, 103, -37, -128, 81, -13, -86, 42, 59, 103, -71, -88, 91, 21, -18, 57, -92, -11, -21, -114, 97, 116, -71, -6, -34, 39, 73, -59, -24, 0, 86, -100, -80, 18, 103, 11, -109, 118, -7, 2, 10, -128, 91, 79, -54, 45, -59, 1, 81, -48, -76, -58, 101, 53, 0, -70, 31, 22, -128, 78, -26, -11, 124, -71, 49, -7, -109, 127, -45, -108, 127, 92, -128, -21, -27, 28, 93, -124, -12, -2, 90, 86, -106, 0, -2, -11, 7, 24, -5, -96, 60, 98, -26, -127, 43, 42, -18, 16, -45, 5, 22, -59, -73, 127, 76, -6, -63, 0, 11, -122, 2, 71, -2, -43, -15, 80, 121, -80, -29, -10, -5, -29, 29, 28, -44, 73, -48, -2, 45, -78, 13, 0, -6, 65, -55, -34, 29, -50, 45, -8, 38, 17, -36, 3, 31, 119, -97, -68, 47, -60, -49, 11, 103, 119, -55, -128, 12, 86, -13, -85, 55, -10, -63, 124, 45, -128, -29, 90, 0, 26, -111, 43, 127, -128, -54, 42, -60, 81, 127, -118, -128, 127, 3, -7, 113, -128, -108, 93, 15, -28, 48, 37, -24, -69, 7, 97, -55, 21, 55, -5, -33, 11, -38, -55, 92, -6, -7, -16, -63, 31, 127, -118, -31, 74, -111, 60, 81, -37, -58, 11, 43, -22, 7, -73, -1, 127, 1, -119, -74, 45, 32, -65, 65, -15, -2, 44, -18, 91, -44, -122, 114, 74, -76, 43, 15, -108, -32, 127, -18, -47, 13, 44, -17, -128, -1, -7, 109, 10, -27, 55, -87, 27, 49, -15, -3, -37, 10, 58, 31, -121, 33, 23, -27, 119, -11, -85, -22, -13, -95, 88, 127, -7, -114, -64, 45, -29, 69, -23, -73, 38, 53, 92, 3, -8, 7, -87, -116, 0, 127, -16, -42, 109, -64, -49, 111, -73, -128, 127, 45, -24, -45, -55, -22, -27, 6, 123, 32, -66, 26, -103, 44, 75, -22, 3, -88, -44, 127, -38, -92, 102, 38, 11, 36, -102, 17, 70, -24, -73, 16, 88, -128, -93, 127, 22, -128, 127, 31, -74, 29, -44, -42, 36, -11, 22, -27, 55, 113, -71, 31, -22, -106, 44, 100, -73, -80, 76, 47, 32, -12, -23, -66, 37, 68, -34, 54, -117, 3, 96, -87, -70, 22, 7, -29, 16, 39, -49, 36, 55, 2, 3, -63, 17, 69, -39, -15, 116, -113, -23, 76, -73, -43, 97, -15, -128, 121, 11, -12, 92, -34, -68, -109, 26, 75, -27, 42, 12, -16, 49, -54, 33, 85, -29, 3, -54, -101, 68, 117, -33, -95, -57, 64, 78, -33, 33, 43, -113, 34, 17, -128, 112, 127, -27, -128, 16, 127, -116, 23, -29, -26, 17, -119, 127, 108, -34, 12, -74, -66, 98, -60, -92, 127, 47, -13, -88, -50, 78, 11, -93, 10, 78, -92, -7, -15, -8, 127, -29, -3, -22, -59, 127, -29, -57, -49, 24, 74, -6, 3, -8, 11, 65, 27, -87, -27, -5, 10, -32, -10, -31, 50, 74, 21, -37, -96, 63, 12, 54, -45, -26, -43, 0, 100, -24, 1, -87, -75, 31, 22, 0, -26, 50, 90, -48, 32, -55, -33, 54, -5, 78, -18, -63, -32, 50, 28, -44, -57, -21, 0, 103, 80, -33, -24, 17, -6, -97, 87, -34, -124, 36, -5, 60, 1, -93, 88, 28, 60, -13, -65, 52, 26, -85, -26, 101, -114, 50, 22, 7, 21, -39, 116, -101, -74, 55, -45, 13, 45, 63, 11, -118, 33, 8, 18, 29, -47, -23, 48, 0, -36, 91, -109, 21, 127, -128, -71, 11, 79, 90, 0, -117, -64, 29, -44, 27, 48, 50, -52, 24, 127, -93, -75, 22, -47, -17, 5, 70, 107, -65, -32, -10, -8, 117, -28, -96, 8, 87, -55, -102, 0, 36, 65, -42, -17, -11, 38, 47, -74, -16, -8, 92, 49, -3, 36, -6, -17, -85, 48, 52, -122, -28, -31, 109, 1, -128, 127, 87, -2, -38, 1, -92, 16, 52, -106, 91, -8, -2, 78, -2, -8, -118, -15, 49, 49, 43, -124, -52, 18, -16, 5, -15, 95, 109, -37, -80, 75, 5, -121, 11, 39, 33, 71, -47, -128, 63, 57, -27, -22, 17, -7, -45, 1, 18, 38, 11, -58, -15, 102, 12, -32, 44, 24, -47, -42, -45, -2, 65, 79, -33, -106, 17, -2, -28, 101, 44, -93, -93, 31, 79, -52, -23, 127, -6, -128, 12, 112, -86, 31, 28, -29, -36, 10, 127, -55, 15, -98, -5, 31, -36, 73, 36, -18, -127, 87, 21, -68, 114, -79, -128, 37, -6, 0, 64, 48, -57, 12, 27, 18, 52, -128, 16, 96, -45, -88, -44, 116, 36, -98, 38, 3, -57, 119, 113, -102, 1, 60, -45, -76, -69, 76, 102, -28, -5, -91, 1, 55, -13, 29, 27, -90, 3, 31, -75, 55, 0, -36, -68, 127, 29, -31, -11, -80, 39, 70, -47, -107, 18, 90, 97, -86, -33, 103, 12, -39, -55, -28, -50, 49, -6, 33, 119, -128, 33, -13, -100, 93, 101, -28, -32, 39, -95, 0, -7, -8, 102, -78, -2, 45, -80, -3, 2, 11, -17, 6, 65, -53, -8, 91, -68, -53, 88, 108, -93, -2, 76, -73, 34, 49, 3, -24, -68, -59, 38, 0, -42, 22, 54, -42, 21, -5, -16, 112, -86, 13, 121, -32, -127, -55, 86, 68, -13, 6, -54, -33, 93, -90, -92, 75, 31, -60, -12, 24, -17, 86, -16, -92, 15, -16, 50, 123, 12, -128, 48, 66, -128, 92, 90, -48, 36, -75, -16, 97, -68, -55, 13, -34, 87, -42, -66, 13, -29, 65, 57, -47, 13, 70, -90, 32, -18, -10, -17, 53, 11, -50, 60, -39, -15, -68, -24, 71, 68, -45, -95, 127, 27, -117, 121, -38, -65, -15, 6, 63, 45, -58, -24, 49, -55, -1, 17, -32, 42, 21, -97, 6, 55, -16, -73, 107, 112, -53, -24, -47, -50, 54, 10, -27, -10, -50, 96, 127, -128, 13, -26, -24, 39, -112, 87, 60, -80, 69, 2, -103, -3, 5, 73, 80, 42, -17, -119, -68, 73, 27, -60, 29, 98, -32, -128, 43, 59, -44, -12, 47, 65, 15, -38, -45, -59, 29, 87, 7, -102, 24, -13, -1, 58, -128, 97, 6, -12, 127, -85, -60, 12, -74, 15, 116, -36, -1, 86, -38, -65, 58, 21, -13, -8, -87, 3, 102, -79, -24, 112, -1, -45, 12, -57, 23, 127, -113, -18, 91, -86, 24, 122, -119, -95, -11, 69, 80, -128, -54, 93, 23, 65, -60, -109, 85, -1, -73, 87, 65, 33, -87, -75, 127, -11, -122, 23, -15, -75, 127, -8, -92, 78, -44, 26, -1, -48, 65, -63, -49, 52, 85, 36, -97, -60, 42, -11, -34, 127, 12, 0, 10, -128, 127, 12, -121, 17, -31, 13, 55, -3, -70, 34, 66, 58, -45, -128, 112, 34, -22, 78, 0, -81, 28, 11, -64, 8, -58, -44, 50, -15, 66, 57, -8, 58, -36, -55, -76, 23, 26, 79, 60, -123, -43, -23, 12, 75, 28, -65, 44, 66, -47, 16, 50, -66, 8, 10, -128, 47, 63, 27, 11, -27, -18, 44, -47, -113, 109, -22, -44, 100, -28, 53, -39, -127, 63, 58, 0, -38, -90, 106, 100, -102, -86, 92, 23, 7, 12, -57, -8, 55, -38, -29, 75, -22, 37, 44, -47, 11, -16, -48, 2, -68, -16, 90, 74, 21, -54, -128, 107, -27, -117, 15, 45, 10, -69, 32, 50, -15, -23, 95, 47, -47, 29, -101, 15, 113, -93, -86, -6, 73, 26, 55, 74, -31, -87, -48, -24, 5, 74, -13, -66, 31, -36, 54, 98, -65, -28, 11, -10, -27, 12, -10, -31, 57, 60, 33, -5, -92, -47, 81, 39, -114, -86, 127, 127, -128, -106, 43, 10, -21, -34, 50, 45, -73, 37, 48, -59, 90, 81, -32, 12, -5, -8, -112, -65, 17, 27, 45, 76, 10, -7, 63, -88, -128, 101, 7, -96, 8, 21, 17, -75, 18, 121, -36, -52, 91, 34, -10, 17, -10, -102, 11, 95, -50, 24, 21, -71, -34, -68, 17, -11, 96, 27, -128, -23, 127, 29, -90, 57, 48, 8, -36, -49, 42, 87, 24, -28, -17, 33, -87, -37, 49, -16, -79, 57, 7, -65, 64, 12, -96, 54, 127, -128, 22, 74, -66, -49, -29, 12, -17, 112, -17, 26, 0, -87, 109, 58, -119, 10, 50, -43, 92, 32, -12, -23, -68, -69, -28, 24, -23, 70, 79, -128, 27, 87, -71, -13, 108, 53, -122, -17, -18, -22, 127, -27, -32, 85, -73, 7, 116, -69, -128, -42, 108, 12, -76, 6, -6, -1, 45, 34, -74, 21, 48, -1, -26, 18, 85, 2, -112, 15, 127, -50, 2, -55, -107, 118, 42, 0, -63, -86, 6, 69, 127, -128, -85, 60, -71, 78, 58, 3, -53, -2, 106, 26, -122, -6, 127, -43, -58, 8, 23, 48, -71, -128, 69, 55, -32, 52, 8, 0, 0, -5, 7, -2, -59, -66, 101, -53, -10, 65, 23, 28, -43, -7, -27, 43, 53, -32, 22, 11, 3, -107, -58, 78, 55, -112, 34, 13, -10, -3, -71, 80, -12, -23, -59, 54, 127, 0, -75, -52, 24, 21, -18, 63, 31, -128, 49, 3, -52, 31, -8, 47, -96, 17, 127, -53, -32, -18, 32, 36, -128, 44, 42, 1, 101, -80, 8, 50, -128, -92, 97, 11, -23, 90, -53, 38, 100, 5, -60, -28, 42, -81, -18, 90, 33, -90, -124, 45, 24, -15, 53, -26, 39, 29, -63, 0, 31, 24, -90, 75, 43, -128, 75, 43, 16, -5, -79, -5, 33, -52, 39, 42, -38, -12, 64, -21, -24, 114, -64, -79, -5, -33, -49, 23, 80, 44, -13, -90, 66, 79, -24, 34, -27, -100, -29, 109, 59, -65, -63, 90, -3, 1, -37, -103, 127, 66, -128, 21, 32, -123, 24, 93, 98, -1, -128, -66, 39, 45, -39, 15, 127, -13, -36, 42, 21, -55, -100, 0, -24, -7, 74, -55, 7, -13, 70, 12, -52, 90, -38, 45, -11, -128, 116, 10, -23, 96, -45, -43, -54, -66, 37, 73, -24, 34, -54, -12, 17, 0, 90, -37, -97, 8, 100, 64, -24, -87, 1, 63, -74, -15, 127, -17, -69, 16, -60, -6, -5, -18, 116, 44, -27, -92, 1, 50, -42, -38, 11, 3, -7, 59, 26, -29, 39, 88, -119, -26, 86, -48, -96, -17, 127, -12, 7, -2, -128, 26, 6, 90, 37, -1, -42, -28, 87, 12, -18, -60, 87, -23, -81, 29, 58, -28, -13, 100, -103, 0, 32, -76, 36, 26, -52, 53, 34, -45, 71, -91, -90, 63, 57, -11, -39, 95, -47, -127, 112, 118, -111, -59, 68, -47, -48, 93, 71, -103, -63, 59, -45, -65, 127, 0, -127, 45, 3, -44, 113, -7, -117, 127, 37, -128, -6, 127, -13, 0, -10, -121, -28, 42, 32, 73, 63, -1, 0, -106, 52, -15, -69, 11, -47, 21, 63, -60, 60, 74, -21, 43, -128, -18, 127, -13, 8, -48, -36, 60, -29, 47, -6, -78, -75, 31, 26, -5, 123, -10, -18, 0, -8, 27, -123, -28, 42, -47, 10, 11, 86, 78, -119, -106, 81, 85, 26, 15, 8, 17, -74, -78, -64, 65, 100, -55, 2, 12, 37, -48, -50, 118, -75, -43, 124, -2, -119, -54, 44, 59, 29, 28, -60, -80, 60, 36, -7, -74, -49, 97, 127, -90, -70, 50, -27, -11, 0, 95, 10, -66, 87, -23, -91, -53, -12, 49, 16, 78, 49, -7, -34, -86, -42, -26, 100, 127, -88, -60, -55, 39, 49, -47, -47, 3, 118, 39, -123, -28, 127, -6, -93, -80, 127, 2, -13, 16, 0, 66, -121, 52, 7, -5, 54, -96, -29, 66, -42, 38, 79, -78, -73, -50, -11, 64, 12, -13, 27, -55, 6, 53, -34, 95, 85, -29, -21, 1, -76, -63, -3, 53, 2, -114, 108, 65, -29, 64, -71, -55, 109, 81, -128, -45, 127, 23, -81, -70, 28, -52, 53, -15, -128, 127, 97, -128, 26, -27, -65, 127, 5, -128, -11, 58, 3, -34, -50, 31, 102, 10, -31, 15, -52, -15, 6, -47, -13, 78, 2, -29, 108, 1, -29, 27, -116, -23, 113, 53, -31, -44, 12, -85, -42, 48, 1, 28, 7, 7, 7, -50, -17, 53, -3, -29, 79, -5, -17, 18, -15, -21, -74, -1, 57, 78, -50, -3, 28, -11, 96, -58, -58, -32, -75, 13, 127, 34, -29, -13, -36, 74, -54, -98, 117, -21, 32, 49, -24, -78, 32, 80, -97, 76, -8, -59, 97, -47, -98, 36, -55, 34, 127, 34, -96, -37, 108, -53, 0, -58, 27, 57, -39, -63, -88, 127, 114, -127, -42, 123, -10, 0, 7, -73, -8, 63, 29, 1, -70, 36, 73, -128, -68, 49, 92, -73, -69, 36, -87, 119, 127, -75, -87, 53, -36, 15, 122, -103, -11, -44, -23, 3, -68, 87, 36, 29, 73, -86, -128, 24, 127, -29, -113, 44, 64, -16, -48, 2, -10, -44, 74, 63, -70, -65, -1, 53, -10, 28, 50, -24, 6, 8, -31, 18, -43, -60, 75, 112, -18, -102, 17, 31, -92, -75, 95, 127, -116, 2, 48, -114, -32, 66, 0, 32, 127, -128, -118, 127, 33, -53, -16, 6, 106, -71, -37, 127, -44, -128, 98, 127, -6, -101, -21, 64, -119, 8, -1, -86, 100, 76, 31, 24, -5, -119, 0, 74, -13, -47, -49, 0, 0, 12, 1, 63, -45, -65, 79, 93, 10, -80, -107, 0, 127, -50, 6, 78, -128, 18, -8, -31, 127, -55, -17, -15, 16, 2, 15, 24, -64, -16, -2, 31, 10, 124, -53, -27, -29, 12, 79, -108, -71, 29, 36, 3, -54, -24, 75, 37, 22, -3, -3, 28, -54, 22, -31, 33, -5, -86, 1, -15, 10, 28, 21, 38, 87, -79, -102, 16, -13, 26, -16, -38, 75, 90, -85, -119, 70, 119, -47, -114, 0, 97, 127, -116, 5, 123, -96, -50, 102, -49, -8, 107, -128, -70, 18, 107, -11, -128, 32, 13, 11, 17, 118, -54, -128, 119, 127, -92, -97, 97, 69, -31, -47, -90, 17, 6, -85, 117, 96, -63, 43, 39, -128, -6, 42, -32, 65, -2, -64, -16, 71, -63, -111, 127, 80, -10, -85, -33, 98, -18, -71, 34, 97, -76, 28, 55, -68, 76, -52, -6, 15, -93, 42, 70, -31, -50, -1, -37, -28, 55, 0, -48, 1, 86, 28, -23, 29, -64, 31, 70, -26, 8, -49, -43, -22, 11, 55, -17, 63, 0, -28, -26, 11, -32, -29, 121, -60, 5, 12, -2, 78, -60, -13, -65, -2, -7, 38, 15, -65, 86, -16, 2, 53, -75, -2, -6, -80, 107, -18, 8, 60, -34, 1, -54, -57, 0, -1, 38, 49, 2, -42, -27, -6, 0, 50, 98, -58, -66, 10, -23, -16, 34, 102, -97, -59, 116, -57, 47, 21, -68, 123, -90, -100, 54, 78, -12, -100, 60, 107, -8, -12, -48, -108, 92, 127, -33, -64, -26, 34, 16, -7, -108, -15, 127, 18, -128, 71, 17, 1, 22, -108, 80, -32, 12, -18, -100, 111, 18, -10, -13, -5, 48, 0, -73, -13, 17, 13, -2, 10, 93, -22, -57, 54, -22, -47, 73, -23, 3, 53, -38, -78, -37, 54, 98, 6, -117, -69, 38, 121, -22, -128, 5, 1, -33, 127, 79, -106, -58, 101, 100, 13, -118, -63, 11, -73, -2, 119, 34, -36, 12, -13, 54, 64, -100, -96, 47, 97, -90, 17, -8, -57, 33, 45, -23, -128, 127, 64, -128, 29, 112, -85, -102, -6, 50, -15, -43, 24, 36, 39, 39, 27, -69, -3, 59, -76, 1, 90, -36, -73, -5, -36, 91, -13, -63, 75, -69, -65, 117, 127, -73, -37, -22, -36, 118, -59, -128, 64, 127, -69, -53, 127, 26, 7, -103, -39, -32, 71, 78, -128, 69, 80, -101, 11, 12, 42, 38, -95, -11, -64, 70, 49, -128, 49, -15, 28, 121, -112, 1, 124, -92, -34, -17, 8, 127, 44, -118, -97, 97, -55, 3, 127, -91, -93, 102, 34, -88, 49, -3, -74, 28, -55, -65, 68, -3, -21, 127, -7, -128, -33, 117, 44, 43, -70, -63, 65, 0, -53, -36, 127, -49, 6, 45, -75, -50, 5, 111, -76, -88, 127, 45, -45, -34, -29, 26, -26, 59, -32, -93, 3, 102, 97, -128, 29, 127, -23, -57, -80, 31, 71, -22, -100, 29, 119, -128, 24, 60, -29, 63, -128, 27, 124, -128, -13, 49, 39, 16, -128, 24, 114, -54, -96, 108, 95, -109, -15, -21, -38, 111, 68, -107, -70, 127, -15, -26, 15, -68, -45, 73, -10, -3, 16, -103, 100, 122, -87, -128, 22, 119, 45, -71, 11, -24, -44, -13, 37, 101, 10, -98, 16, 123, -42, -31, -43, 58, -69, -101, 70, -43, -39, 97, 53, -36, -37, -29, 47, 28, -71, 11, -2, 70, -2, -121, -3, 112, 127, -106, -59, 64, 70, -58, -128, 34, 98, 49, -34, 12, -39, -50, 107, 3, -91, -80, 58, 80, -33, -22, -37, -74, 52, 127, -60, 18, 18, -57, 114, -54, -98, 43, 93, 13, -128, 17, -18, 17, 97, -34, -70, -76, 65, -22, 95, -23, -33, 32, -97, -2, 73, 8, -68, 71, 49, -79, -10, 32, 74, 3, -124, -5, 21, -39, 117, 57, -128, 69, 91, -107, -6, 47, -128, 70, 127, -119, -60, 0, 60, -28, -50, 121, -70, -42, 44, 43, 17, -127, 39, 10, -66, 86, -21, 18, 81, 31, -52, -47, 73, -65, 0, -27, -57, 86, -24, -8, -55, 22, 127, -38, -75, 38, 5, -15, 43, 1, -101, 42, -2, 36, -6, -128, 107, 18, -7, 111, -106, -86, 57, 12, 80, 1, -128, 91, -34, -54, 86, 31, 18, -128, 48, 37, 21, -52, -73, 96, -48, 1, 42, -27, 2, 47, -55, 31, 78, -109, -70, 96, 13, -97, -49, 124, 66, -33, -55, -54, 127, -44, -95, 45, -42, 43, 13, 27, 86, -121, -107, -11, 127, 96, -49, -27, -76, -49, 87, 10, -28, 3, -39, -15, 85, -24, -76, 127, 50, -13, -52, -42, 116, -24, 2, -34, -106, 11, 75, -16, -55, 108, -42, -17, 39, 22, 79, -54, -92, -11, 31, 71, 69, -42, -23, 66, -85, -68, -16, 13, 64, -31, -52, 21, -32, -48, 127, -48, -106, 12, 97, 44, -28, 69, -65, -24, -49, 27, 11, 11, 5, -106, 101, -24, -38, 112, 32, -50, -2, 42, 5, 17, -32, -98, 27, -42, 44, 80, -101, 43, 5, 36, 10, -79, -24, 54, -59, -28, 18, 27, 6, 24, -10, -66, 48, -78, 68, 21, -63, 127, -18, -128, 111, -1, -43, 88, -93, 29, 108, -18, -73, -36, 28, 80, 6, -70, -63, -32, 85, 107, 2, -128, -44, 69, 49, -44, 0, 34, 18, 48, -128, -66, 98, -2, -88, 90, 80, -2, -88, 28, -26, -34, 88, -117, 0, 57, 2, -43, 87, 43, -37, -2, -37, 74, -39, -107, -26, -13, 75, 38, 64, -47, -27, 26, 0, -32, -93, 31, -6, 17, 117, 78, -128, 29, 13, -70, 54, -52, -31, 33, 63, -60, 50, 32, -117, 1, 39, -8, 49, -31, 22, -26, -17, 0, -2, 119, -55, -22, -7, 55, 5, -109, 6, -21, 75, 100, -74, -27, -38, -66, 80, 75, -47, 10, -43, 48, 127, -112, -37, 98, -16, -18, 1, -58, -38, 102, -12, -33, 58, -100, 49, 45, -128, 92, 18, -128, 34, 102, 28, 0, 42, -128, -49, 11, -66, 101, 64, -42, 66, -49, -42, 59, -6, 0, 28, -57, -100, 1, 71, 38, -55, 54, -34, 16, 102, -128, 0, 12, -85, 127, 109, -118, -112, 43, 11, 10, 49, 38, -13, -102, 27, 28, 69, 81, -128, 36, 29, -71, 54, 18, 70, -79, -107, -34, 87, 26, -87, 24, 59, -50, -29, 33, 86, 112, -128, -93, 117, -47, 18, 127, -128, -39, 11, -50, 92, -23, 38, 101, -55, -107, 64, -22, -128, 17, 88, 127, -96, -128, 54, 109, 59, -59, -3, 42, 12, -95, -121, 24, -10, 113, 10, 0, 26, -127, 88, 27, -15, 95, -3, -79, 17, -64, 0, 121, -117, -97, 8, 98, -10, 23, 113, 0, -113, 10, -15, -73, 28, 31, 21, -28, 96, -87, -27, 95, -37, 42, 70, -101, -128, 79, 49, -27, 2, -63, -59, 39, 100, -55, -36, 111, 6, 18, -10, 7, 90, -128, -39, 70, -100, 88, 64, -128, 69, 31, -128, 11, 63, -79, 65, 73, -128, 22, 91, -22, -47, -79, 112, 127, -128, -18, 103, -11, -102, 39, 107, 12, 10, -90, -5, -47, -58, 1, -37, 42, -24, 80, 74, -114, -22, 6, -64, 127, 24, -75, 22, 23, 18, -59, -21, 1, -29, 24, 116, -60, -47, 18, 33, 103, 12, -74, -95, -21, 116, 76, -36, -57, 17, 74, -55, -103, 26, 11, -23, -18, -69, 127, 26, -98, 59, 75, -80, 15, 11, -100, 36, 16, 15, -17, 59, -1, -81, 49, 22, -52, -10, 50, -6, -31, -29, 87, 113, -42, -128, 17, 69, -74, 39, 3, -97, 80, -34, -24, 127, 38, -100, -75, 39, 78, 42, -128, -100, 65, -22, 74, 114, -85, -64, -2, -15, 0, -28, -2, 5, 42, -17, 63, 59, -74, 87, -60, -128, 13, 102, -2, -102, 6, 13, 42, 112, -17, -98, -29, -27, 17, 85, 7, 3, -13, -22, -44, -8, -1, -59, 18, 95, 15, -31, -8, -43, 122, 108, -101, -81, -7, 8, 44, 37, 11, 12, -114, -10, 96, -80, 13, 91, -21, 15, 38, -78, 29, 69, -128, 34, 65, -128, 7, 55, 0, 54, 44, -128, 34, 87, 16, -70, -128, 97, 108, -98, -60, 121, 23, -18, -38, 7, -38, -21, 6, 21, 109, 16, 1, -116, -29, 127, -95, -123, 75, 114, -24, -128, 64, 102, -10, -44, 31, 49, -69, 44, -50, -8, 81, -66, 66, -78, -26, -10, -12, 59, 12, 66, -100, -39, -22, 80, -1, -128, 127, 58, -39, 27, -97, 32, 88, -103, 38, 60, -18, -100, -12, 127, -68, -36, -28, 17, 17, 5, -13, -13, 66, -103, 65, 48, -8, -43, -21, -7, -79, 10, 10, 64, 101, -92, -102, 116, 17, -43, 13, 21, 76, -108, 26, 66, -112, -15, 39, -26, -34, 43, -11, 32, 97, -70, -107, 117, 64, -23, -39, -90, -34, 45, 127, 1, -70, 5, -7, -32, -50, -42, 127, 17, -95, 27, 34, 92, -47, -32, -42, -59, 127, 64, -128, 39, -2, -69, 33, 17, 73, -7, 23, -17, -93, 60, 26, -128, -38, 117, 80, -88, -69, -28, -27, 3, 66, 11, -49, 42, -17, -5, 103, -36, -39, 111, -71, -88, 55, 81, -33, 15, 85, -128, -101, 0, 127, 127, -117, -73, 123, 5, -2, 2, -76, 63, -50, -117, 106, 15, -109, -18, 11, 123, 85, -69, -34, -75, 18, 81, -53, 42, 33, -86, 24, 75, 31, -27, -49, -18, 66, 27, -124, -98, 73, 80, 45, 54, -97, -55, 18, 13, -8, -47, 90, 81, -87, -124, -7, 127, -6, -107, 98, -34, -119, 127, 47, -70, -3, -7, 1, 16, 57, 6, -116, -2, 34, -86, 55, 55, 23, 34, -128, 50, 5, -10, 60, -108, -44, 22, 28, 66, 3, -50, 43, 2, 2, 52, -112, 15, 111, -112, -54, 17, 78, 33, -112, 53, -8, -34, 127, -121, -80, 34, 28, 81, 10, -31, -91, 10, 81, -16, 28, -34, -49, 78, -36, -45, 59, -90, 38, 124, -52, -112, 13, 127, 0, -48, -28, -36, 54, 39, -47, 58, 31, -29, -91, -81, 80, 55, 27, 2, -42, -85, -87, 6, 127, 93, -109, -52, 112, 103, -108, -8, -37, -68, 38, 26, -17, 49, -3, -65, 121, -66, -5, 3, 5, 98, -28, -128, 18, 127, -33, -31, 44, -50, -106, 49, 45, -100, 75, 93, -10, -1, -12, 36, -24, -23, -57, -45, 18, 88, -17, -108, 42, 0, -17, 10, 28, -44, -1, 112, 10, -128, 66, 36, -76, 33, 63, -5, -128, 108, 71, -48, 22, 42, -44, -109, -31, -37, 69, 26, 12, 102, -2, -42, -93, -66, 127, 108, -68, -128, 74, 27, -37, -7, 29, 2, -76, 103, 24, -26, -16, 28, -54, -101, 107, 15, -64, 95, 39, -128, 17, 103, -45, 55, -8, -34, -53, -15, -10, -31, 42, -18, 15, -48, 79, 127, -117, 0, 54, -100, -27, 74, 60, -100, -107, 97, 127, -54, -87, 73, 36, -75, 38, 108, -33, -128, -38, 109, -66, 1, 97, -39, -53, -22, 11, -6, 100, -42, -90, 106, -13, -74, 101, 68, -59, -43, -39, -73, 119, 103, -117, 68, -29, -87, 11, 10, -11, 34, 127, -127, -73, 3, 74, 86, -119, 49, -2, 23, -12, -90, 50, -69, 76, -23, -2, 8, -58, 12, -10, 92, -1, -63, -12, -45, 100, 33, -96, 102, 53, -128, -12, 49, 23, 0, -76, 116, 16, -128, 49, 3, 10, 69, -64, -5, 22, 0, 64, -39, -36, -2, -15, 88, -42, 12, 28, -48, -71, 64, 73, -128, 3, 29, -11, -3, -80, 127, 17, -112, -8, 93, 90, 5, -37, 6, -57, -59, 64, -50, -34, 60, 124, -3, -123, 13, 119, -6, -71, 26, 45, -107, 18, 47, 15, -48, -38, -5, -108, 101, 123, -6, -128, 5, 18, -26, 81, -86, 18, 57, -47, 5, 68, -50, -106, 66, 64, 2, -63, -52, 38, 26, -1, -12, -43, 26, 113, -45, -23, 96, -65, -2, -49, -93, 70, 45, 2, 7, 38, -21, 28, -18, -128, 48, 123, -33, -60, -53, 2, -12, 68, 1, -13, 127, -58, -112, -49, 31, 54, 45, 5, -95, 37, 101, -91, 54, 45, -128, 18, 52, -90, 118, 0, -128, 42, 78, 44, -69, 59, 11, -87, 78, 34, -102, 45, 106, -24, -36, -57, 76, -6, -97, 36, 103, -98, -96, 111, -29, -15, 65, 53, -80, 1, 26, -18, -31, 27, -24, 0, 11, -86, 58, -47, 68, -22, -78, 127, 0, 7, 11, -65, -24, 43, 26, -6, -49, 12, 66, 3, 32, -78, -88, -13, 18, 26, 1, 29, 17, -21, 13, -63, 17, 24, 17, 58, -15, -29, -85, 36, -13, -76, 114, 111, 21, -96, -69, 102, 32, -50, -43, -65, -27, 0, 127, 127, -66, -123, -75, 18, 13, 31, 21, 79, -1, 2, 34, -50, -98, 58, 68, -128, 76, 96, -74, -48, -42, 49, 113, -38, 29, 11, -128, 98, 18, -98, -6, -32, 54, -5, 0, 43, -10, -59, -32, 86, -47, 15, 86, -113, 26, 65, -2, 21, 36, 33, -48, -114, -81, 127, -13, -10, 38, -76, 58, -1, -65, 12, 75, -16, 7, 66, -47, -80, 23, 12, 8, 29, -12, 27, -81, -95, 70, 18, 78, 27, -31, -73, -22, 50, 21, 44, 3, -69, 0, 116, -8, -103, 47, 11, -128, 90, 69, -42, 31, -33, -1, -13, 60, -23, -12, 28, -70, 12, 66, 54, -37, -118, 36, 23, -36, 2, 10, 11, -66, 36, -29, 64, 127, -128, -10, 121, 1, -79, -81, 91, -63, -52, 127, -59, -85, 8, 87, 32, -58, -53, -66, 127, 0, -98, 15, -48, 97, 112, -81, 11, 6, -116, 39, 26, -27, 107, -23, -127, -3, -23, 127, -12, -15, 116, -90, -109, 49, 97, 22, -57, -57, 90, 70, -101, -101, -1, -45, 121, 86, -49, -100, 81, 1, -78, 85, 15, 22, -74, -27, 117, 7, -16, -3, -117, 55, 22, -76, 66, -53, 28, 111, -47, -29, 59, 38, -32, 13, -33, -119, 31, 66, -85, 57, 103, -39, 0, -90, -95, 60, 57, 38, 37, -23, -128, 29, 127, -92, -29, 50, -109, -1, 127, 24, -79, 44, -18, -91, 49, 98, -36, 8, -47, -29, 107, -123, -58, 80, -11, 66, -17, -95, 26, -49, -3, 15, 108, 70, 10, -95, -124, 95, 92, -97, 8, 71, -37, -12, -34, -18, 32, 107, 12, -22, -2, 26, -108, -92, 11, 16, 117, 70, 3, -128, -10, 48, -36, -6, 44, 32, 21, 58, -78, -60, 0, 85, -18, -128, 17, 127, -55, -60, 3, 15, 54, -86, 55, 124, -69, -58, -45, 65, 33, 1, -28, -3, 81, -50, -92, -36, 127, -2, -128, 42, 127, -31, -52, 57, -3, 33, -57, -12, 91, -128, 7, 127, -109, -12, 8, -58, 91, 43, -18, -37, -32, -15, 49, -32, -90, 11, 90, 57, 21, -65, -88, 124, -80, 6, 68, -128, 112, 103, -57, -95, -88, 127, 103, -17, -17, -123, 43, 6, 11, -21, -10, 109, -32, -6, -53, -26, 0, 13, 48, -12, -32, 1, 12, 55, -45, -1, 27, -15, 17, -3, -55, 38, 103, -60, -69, -31, 96, -49, -13, 22, -112, 81, 3, -48, -23, 64, 58, -90, 76, 52, -58, 1, -68, -75, 127, 47, -128, 127, 8, -128, 127, 70, -128, -27, 55, -37, -26, 37, 64, 100, 32, -87, -23, -42, -74, 0, 65, 74, -90, 43, 119, -12, -27, -1, -121, 21, 127, -124, -106, 101, 43, -66, 32, -28, -50, 24, 68, -15, -102, -3, 88, -1, -24, 1, -91, 55, 127, 10, -85, -29, 12, -6, 12, 96, -38, -18, -6, -64, 16, 96, -42, -86, 98, 33, -86, -43, 68, -50, -66, 29, 75, 69, 2, -128, 36, 127, -119, -102, 76, -17, 44, 74, -29, -45, 2, 101, -24, -28, -7, -91, 16, 122, -37, 18, -37, -113, 79, -42, -69, 48, 109, -50, -76, 127, -58, -107, 95, 96, -43, -49, -73, 10, 127, 11, -33, 8, -59, -128, 59, 52, -54, -13, 10, -2, 75, 71, -128, 54, 15, -44, -2, -23, 103, -97, -92, 23, 29, 114, 93, -48, 1, -75, 5, 44, -8, -75, -3, 32, -93, 32, 100, 5, -95, -22, -27, 7, 69, 85, -3, -49, 8, -39, -70, 58, 88, 65, -96, -124, 39, -39, 111, 39, -124, -15, 79, 36, 18, 38, -91, -100, 107, 121, -128, -54, 15, 60, -11, 31, 113, -128, 10, 36, -49, 58, -28, -10, 66, -85, 18, 127, -100, -23, 57, -22, -12, -75, -80, 127, 119, -16, -57, -1, -17, 2, 43, 10, -24, -43, -28, -23, 15, 32, -57, 36, 127, -128, -93, 73, 10, -13, 64, -53, -75, 8, 79, -11, -47, 33, -58, -3, 12, 64, 50, -78, 32, 122, -122, -119, 127, 16, -36, 76, -97, -42, 50, -24, 69, 39, -128, 49, 127, -64, -50, -76, 76, 28, -65, -6, -48, 97, -15, -12, 63, -1, -75, 27, 58, -121, -18, 127, 32, -74, -16, 7, 31, 2, 2, 0, -48, -50, 116, -16, -12, 98, -128, 13, -8, -112, 88, 98, -26, -87, -31, -7, 93, 50, -53, -12, 31, -45, -37, 92, -48, -23, 97, -22, 39, -7, -128, 81, 96, -33, 37, -11, -36, 31, -59, 6, -18, -90, -12, 127, -7, -128, 11, 18, -12, 45, 127, -53, -97, -5, -39, 127, 31, -128, 81, 66, -24, 65, -70, -116, 27, 88, 31, -10, 37, -50, -128, 119, -2, -85, 48, -15, -12, 27, 15, -15, -49, 39, 127, -11, -91, -11, 38, 37, -60, -68, 68, 54, 68, -59, -88, 33, -15, -64, -16, 59, 127, -57, -16, 38, -31, 5, 5, -29, -74, 66, -31, 58, -29, -16, 109, -87, 43, 5, -127, 37, -7, 55, 74, -128, 65, 116, -101, -128, 34, 97, -18, -69, 15, 90, 71, -106, -59, 8, -58, 15, -2, 65, 66, -118, 55, 53, -65, 60, 18, -68, 31, -6, -55, 121, -3, -122, -27, 103, 78, -88, 1, 31, -118, 75, 75, -128, 39, 18, -68, 111, 44, -45, 55, -90, -34, 95, 17, 54, -128, -31, 54, -23, 91, -36, -91, -21, -44, 106, 127, -128, -55, 127, -90, -64, 127, 60, -109, -70, 22, -23, -17, 58, 113, -96, -128, 74, 127, 12, -17, 43, -100, -123, 42, 98, 10, -92, 64, 81, 8, -64, -59, 95, -71, -54, 73, -54, -52, 107, 32, -103, 8, 38, -1, 92, -2, -128, 42, -1, -10, 124, -55, 11, 36, -76, -63, 78, 32, -85, -16, -57, 97, -12, 5, 114, -86, 23, 44, -65, -106, -3, 59, 39, 102, -127, -16, 92, -78, 68, -60, -38, -10, 21, 101, -58, -78, 43, 113, 37, -118, -44, 112, -27, -88, -55, 70, 48, 48, -66, -64, 49, 3, -31, -10, 43, -87, 79, 127, -123, 13, 75, 11, -57, -29, 100, -44, 11, -64, -111, -5, 63, 113, 1, -16, -26, -54, 63, -34, -98, 11, -13, 92, 42, -39, -15, 15, 27, -74, -2, 63, -57, 75, 112, -128, -88, 127, 73, -81, -92, -5, 127, -86, -8, 127, -128, -66, 32, -44, 55, 59, 7, 1, -52, 2, -34, 59, 100, -45, 16, -85, 8, -8, -49, 74, -57, 91, 2, 10, 0, -54, 100, -119, 44, 27, -128, 127, 48, -128, 52, 13, -124, 16, 59, 58, 22, 68, -114, -24, 98, 12, -15, 3, 22, -33, -24, 29, 23, -59, -32, 47, 54, -21, -58, -31, -1, 3, 8, -2, 69, -60, -8, 95, -22, 6, -42, -66, -27, -12, -7, 69, 91, -5, -64, 34, 119, -128, 0, 86, -17, 55, -66, -26, -70, 54, 68, -8, -38, -95, -1, 69, 103, -109, 22, 113, -13, 2, -121, 12, 7, -71, 38, -32, 1, 90, 81, -100, -127, 87, 15, -24, 111, 8, -106, 43, 29, -128, 17, 47, -48, 64, -38, -23, 100, 23, -36, 49, -31, -24, 0, 27, 8, -121, 101, 37, -90, -70, 73, 48, 32, -26, -128, 103, 119, -93, -2, 39, -106, -65, 101, 12, 58, -32, -26, 123, -113, -75, 49, 60, -39, -43, -22, 95, 2, -76, 64, -68, -16, 106, -13, 17, 0, -109, 95, 21, -128, -2, 127, -5, -76, 76, -24, -5, -23, -86, 119, -21, -128, 6, 18, 127, -8, -11, 38, -32, 54, -71, 0, 98, -107, -11, 111, -63, -79, -12, 66, -21, -37, 95, -59, -108, 45, 54, -5, -33, 50, 39, 21, -44, -111, -10, 95, 91, -44, 2, 50, -79, -60, 17, -34, 57, 21, -63, 53, 79, -42, -49, -37, 88, 97, -49, -54, -58, 103, -31, -57, 49, 43, -2, -113, 36, -31, -66, 100, 28, 0, 52, -86, -74, 119, 45, -54, 29, 68, -92, -18, 65, -128, 68, 127, -128, 16, 64, 15, -50, -78, 90, 64, 21, -74, -70, -65, 78, 39, -118, -12, -5, 42, 103, 10, -109, -36, 127, 27, -68, 21, -8, -93, 57, 127, -42, -93, -57, -21, 93, 86, -11, -109, -15, 119, 53, -42, -58, -32, -43, -5, -15, -23, 57, 0, -37, 78, -55, 63, 127, -106, -31, -49, -36, 101, 54, -10, 5, -48, 7, 58, -128, 55, 127, -91, 44, -44, -118, 127, -23, -52, -1, -26, 124, -6, -45, -54, -59, 45, 37, 68, 10, -73, -53, 48, 80, 28, 7, -74, 5, 57, -18, -81, -8, 127, -63, -81, -48, 91, 24, -80, 102, 34, -26, -112, 36, 88, -21, -3, 22, -2, -88, -76, 93, 92, -79, -32, -57, 78, -8, -6, 91, -86, -54, -42, 73, 39, 38, -33, 21, 17, -37, -34, 1, 127, -54, -71, 38, -39, -33, 28, 54, 81, -81, -86, 101, -17, -97, -3, 44, 66, 1, 2, 54, -45, -52, 17, -52, -26, 68, -60, -63, 127, -54, 1, 1, 12, -8, -6, 127, -117, -70, 127, -66, -57, 123, -12, 31, -45, -76, -5, 55, 59, -15, 28, -39, -16, 16, -80, -2, 95, -60, -98, 92, 55, 21, 42, -128, -12, 68, -63, -36, 74, -23, -48, 17, -6, 88, -69, 16, 122, -73, 23, 74, -121, -86, 74, 73, 43, -111, -63, 103, -2, -15, 57, -50, -28, 13, -43, -6, 102, 18, -44, -29, 24, 22, 3, 74, -24, 0, -31, -128, -45, -1, 116, 63, -128, 69, -1, 5, -2, -52, 48, 28, -15, -59, 121, 59, 6, -69, -64, 75, 0, 5, -6, -93, -28, 100, 91, -63, -5, 23, -119, -64, 0, 127, 96, -128, -59, 127, 52, -101, -101, 29, 27, -12, -32, 100, 6, -127, 63, -39, 75, 127, -73, -109, -37, -18, 124, -3, -64, 127, -93, -113, 127, 13, -59, 101, 31, -128, -1, 127, -128, -128, 75, 71, -28, 74, -17, 3, -2, -128, 59, 26, -66, 96, 49, -31, 5, 50, 58, -3, -32, -85, -11, -28, 58, 119, -28, -128, -5, 102, -15, -92, -86, 95, 81, -29, -12, -48, 55, 39, -65, 45, -49, -31, 127, 5, -91, -1, 7, 55, 42, -128, 22, 42, -116, 80, 75, -112, 12, 55, 26, 68, -121, 23, 95, -22, -85, 15, -18, -69, 118, 55, -88, -91, 117, -54, -102, 38, 28, 5, -58, 11, 92, 38, -96, -54, 127, -17, -63, 27, 49, 68, -17, -59, -39, 86, 55, -64, -69, 60, -12, -8, 45, 33, -116, -43, 127, -74, -128, 45, 91, 28, -47, 23, 63, -91, -7, 81, -90, 6, 15, -128, 108, 127, -123, -81, 55, 12, 70, 0, -87, 3, -22, -3, -5, 44, 123, -17, -128, -47, -5, 100, 11, -22, 119, -65, -102, -3, 57, 87, -108, -60, 117, -78, 45, 127, -128, -6, 127, -58, -22, -50, -81, 36, 64, 85, 0, -37, 65, -97, -106, 60, 75, 59, -112, -128, 59, 113, -23, -38, 88, 75, -128, -93, 15, -28, 127, -18, -69, 95, 42, -106, 49, 79, -128, -13, 5, -58, 7, 113, 0, -39, 12, -3, 39, -22, 48, 59, -70, -108, 49, 127, -26, -74, -57, -70, 114, 68, -38, 59, -93, -119, 11, -13, 116, 121, -23, -80, -23, -42, -5, 127, -33, -88, 49, 0, 64, -24, -28, 0, -109, -17, -16, 117, 127, -7, -128, 22, 113, -47, -37, -10, 3, 0, -11, -31, -7, -65, 96, 75, -59, -1, -32, 2, 5, 64, -65, -13, 93, -103, 26, 78, -92, -53, 79, 75, 44, -68, -79, 6, -12, -24, -50, 18, 76, 76, -31, -109, 17, 16, -6, 75, 63, 22, -113, -121, 26, 3, -15, 87, 103, -86, 26, 27, 0, -75, -47, 127, -127, 17, 98, -128, 52, 29, 2, 28, -52, 68, 39, 3, -86, 10, 66, -78, -8, -2, 2, 0, -79, 45, 102, -13, -90, 10, 97, -11, -109, 16, 64, -107, 69, 24, -128, 0, 127, -21, -128, 102, 45, -50, 73, 54, -10, 13, -128, -7, 118, -22, -98, 49, 100, 6, -57, -59, 79, 7, -47, -36, -11, 10, 32, -2, 8, 75, -2, -74, 0, -11, -37, 31, -11, 48, 42, -90, 38, -3, -36, 27, -53, -49, 109, -5, -128, 74, 52, -70, 73, 68, -128, 81, -12, -76, 127, -97, -50, 71, -121, 57, 107, -107, 18, 12, 52, -27, -111, 127, -17, 0, 58, -55, -78, -34, 127, -69, -97, 127, -48, -70, -7, -52, 7, 37, 80, 2, -79, 79, -12, -117, 127, -43, -3, 127, -128, -23, 116, -108, -10, 102, -66, -87, 102, -24, -48, 113, -2, -100, -47, 127, 50, -44, 34, -49, -64, 11, 90, -76, -128, 102, 106, 43, -111, -93, 32, -13, 0, 75, -22, 32, 75, -18, 6, -55, 53, -15, -123, 81, 47, 1, 76, -123, -24, 11, -108, 95, -2, -43, 78, -18, -65, 103, 7, -102, 15, 27, 90, -37, -33, 2, -12, -38, 6, -12, 3, 127, 1, -90, -44, 26, 81, 66, -34, -81, -97, -23, 106, 108, -32, -128, 27, 78, -88, 44, -23, 47, 7, -50, 5, -49, 6, -49, 43, 63, 78, 42, -128, -74, 107, 81, -93, -101, 71, -3, -43, -6, 90, -33, 21, 100, -39, -37, -65, 31, 13, 66, -17, -5, 48, -17, -53, -8, 17, -86, -44, 127, -31, -13, 45, -45, -16, 39, 100, -128, 31, 47, -60, 121, -27, -64, 63, -22, -57, -11, -43, -36, -6, 64, 44, -74, 43, 119, -68, -100, -10, 75, 69, 13, 0, -109, 39, 119, -106, -63, 1, -70, 127, 101, -80, -18, 53, 23, -122, -37, 58, 31, 42, -71, 10, 0, 32, -28, -39, 127, -69, 27, -26, -57, 29, 27, 57, -57, -52, -50, 0, 52, 52, -10, -69, 24, 64, 48, -11, -16, -65, -38, 60, 42, -24, -92, 65, -36, -36, 27, -69, 71, 29, -85, 101, 57, -128, -63, 114, 122, -124, -70, 22, -45, 60, 29, 26, -38, -1, 17, 10, 16, -38, 116, -85, -49, 93, -85, 11, 112, -44, -57, 0, 78, -10, -17, 12, -90, 63, 15, 22, 23, -88, -11, 34, -48, 63, 3, -42, 92, -101, -103, 60, -3, 73, -13, -34, 36, 39, 24, -38, -29, -106, 59, 75, -26, -12, 18, -75, 34, 28, -121, 127, 92, -26, 10, -98, -64, 53, 108, 58, -119, -95, 88, -37, -80, 127, 75, -70, -68, -2, -18, 0, 127, -71, -128, 127, 85, 15, -117, 16, 53, -71, -24, 70, 21, -92, 18, -13, 92, -52, -22, 122, -87, -68, -12, 26, 100, -65, -38, 60, -28, -49, -2, 16, 101, 16, 3, -55, -109, 91, 0, -10, -34, -7, 37, -34, 52, 76, 17, -78, 11, 18, -59, -15, -10, -1, 5, -29, 71, 18, -64, -54, 100, 38, -34, 45, -59, 38, 55, 27, -121, -106, 32, 22, -2, 108, -5, -123, 0, 102, 3, -128, 127, 16, -29, 111, -36, -90, -100, 39, 10, 88, 26, -15, -10, -128, 74, -21, 32, 43, -85, 28, 107, -44, -2, 26, -38, 54, 12, 10, -63, -60, 36, 92, -63, -39, 100, -50, -91, 111, 10, -76, 66, 7, -47, -32, 0, 98, -38, -65, 74, -88, -43, 127, -37, -87, 3, 10, 70, -53, 28, -2, -10, -1, -93, 113, 27, -102, 100, -26, -101, 73, -18, -59, 27, 43, 48, -16, 6, 100, -111, -88, 123, 45, -16, 0, -85, -86, 69, 74, 38, -59, 2, 3, -122, -31, 97, 127, -55, -91, 15, -32, 68, 87, -102, 0, -17, 58, 47, -18, 32, -33, -106, -71, 127, 119, -96, 18, -48, -59, 127, -60, -92, -28, 86, 2, -93, 1, 96, 53, -2, 43, -73, 16, -50, -92, 127, -32, -48, 119, 11, -69, -60, -7, 66, -39, -8, 44, -128, 93, 69, -7, -80, 6, 79, -100, 1, -18, -53, -13, 122, 39, -103, -11, 80, 65, -33, 58, -90, -113, 127, 66, -66, 7, -102, 0, 106, -58, -76, 79, 22, -15, 0, -27, -31, 33, 127, -128, -2, 103, -128, 3, 34, 17, -5, -26, 106, -117, -57, 111, 1, -66, 1, -37, 58, 123, -128, -112, 42, 73, 70, -79, -70, 26, 42, 33, 0, -52, -68, -2, 119, 116, -11, -78, -106, 44, 45, -57, 17, 36, 63, -68, 27, 0, -92, 64, -36, 16, 12, 45, 38, -90, -7, 50, 54, -24, -24, 73, -79, 22, 8, -122, 74, 11, -106, 37, 17, -79, 108, 127, -68, -123, 22, 114, -73, -128, 101, 111, -23, -96, 38, 81, -36, 21, -114, -3, 116, -36, 34, 42, 8, -81, -95, 16, 26, 73, -23, -53, 29, 48, 27, 0, 28, -111, -119, 127, 23, -12, 27, -96, 17, 44, -22, 45, -86, 22, 127, -33, -43, 0, -36, 17, -34, 0, 45, -128, 13, 37, -18, 101, 10, -57, 58, 34, -96, -13, -34, 0, 34, -38, 95, 43, -38, -13, -79, 26, 127, -38, -60, 78, 1, -63, -78, -31, 2, 8, 74, 7, 10, 0, -81, 36, 12, -6, -10, -90, 1, 88, -21, 26, 1, 18, 44, -128, 13, 60, 95, 5, -121, 21, 88, 8, -42, -96, 11, 118, 27, -98, -75, 0, 57, -21, -29, 64, -16, 15, -45, 58, 29, -16, 73, -109, 15, 48, -128, 73, 127, -45, 8, -58, -33, 55, -39, 11, -24, -96, 3, 124, 43, -15, 37, 2, -29, -93, -38, 93, 47, -52, -112, 59, 91, 6, -2, -68, -8, -21, 3, 78, 3, -78, 49, -64, -21, 127, -66, -106, 3, 65, 63, 29, -102, 3, 113, -29, -28, 2, -90, -1, 22, -32, -8, 32, 18, 13, 26, -111, 10, 1, -12, -10, 13, 111, -6, -98, -5, 111, 48, -102, -109, 6, 98, 5, -24, -10, -50, 70, 119, -49, -50, -55, -27, 92, -68, -44, 43, 45, -2, -54, 55, 34, -55, 27, -28, -73, 15, 127, -43, -5, 127, -128, -128, 49, 85, -12, 54, -28, -128, 127, 91, -23, -55, -11, 6, 29, -15, -73, 42, -26, 6, 93, -5, -59, 55, 55, -8, -53, -78, -65, -18, 127, 27, -88, 52, 107, -128, -22, 34, -117, 26, 59, 80, 38, 22, -109, 15, -22, -73, 73, 43, -55, -127, 103, 18, -97, 12, 127, -26, 5, 27, -128, 109, 127, -45, -103, 28, 44, -55, -50, 60, 96, -122, -16, 66, -54, -28, 65, -50, -70, 123, 53, -80, -24, -26, 101, -28, -26, 127, -108, -50, -15, 17, 127, -93, -13, 90, -15, -1, -70, 3, 36, -92, -57, 3, 36, -1, 96, 21, -13, 34, -17, 27, -112, -86, 1, 3, 127, 80, 7, -78, -18, 13, -73, 29, 50, -63, 8, -16, -34, 11, -48, 76, -21, -42, -22, 119, 114, -17, -6, -107, 17, 91, -21, -85, -85, 93, 64, -68, -13, 0, -48, 93, 109, -55, -2, -66, 2, 113, -54, -128, 63, 23, -65, 39, 3, 5, -8, 8, 48, -93, -74, 122, 98, -13, -128, 34, 50, -10, 76, -10, 3, 21, 3, -128, 39, 50, -76, -37, 23, 15, -87, 118, 75, -98, 12, 97, 7, -52, 0, 0, -49, 55, 17, -85, -59, 44, 29, 55, -63, -60, 58, 18, 85, 10, -128, 7, 90, 8, -74, -98, 11, 106, 42, -128, 76, 1, -81, 29, -31, 63, 39, 28, 60, -36, -3, -16, -96, 8, 88, -68, -29, -6, 13, 57, -6, -28, -81, 43, 39, 47, 8, -22, 6, -8, -21, -48, 28, 10, 65, 22, -119, 2, 118, 5, -128, -57, 90, -42, -33, 17, -34, 38, 124, -36, -24, 27, -112, -12, 1, 31, -13, 87, 54, -128, 91, -2, 17, 57, -128, 10, 27, -31, 103, 17, -18, 7, -21, -49, -79, 39, 27, -38, -27, 32, -22, 13, 0, -42, 102, 32, -81, 64, 0, 50, 11, -123, 5, 7, 73, 42, 29, -58, -116, 48, 127, -71, -128, 127, 109, -128, -74, 100, 42, -96, -74, 118, 127, 2, -21, -47, -16, -34, -50, 93, -33, -106, 7, 11, 65, 36, 28, -63, -85, 39, 0, -17, 48, 88, -21, -101, -23, 114, 18, -39, -68, 12, 44, 36, -43, -39, 64, -8, 39, -66, -36, 91, 81, -122, 3, 111, -128, 13, 81, 6, -36, -60, 58, -88, -50, 102, -31, 37, 18, -85, 66, 78, 1, -128, 22, 49, -53, -52, 21, -8, 65, 18, -24, 55, -66, 57, -66, -98, 122, 107, -103, -79, -17, 81, 127, -114, -66, 49, -18, 45, 88, -38, -86, 29, -57, -74, 0, 92, 121, 27, -123, -111, 109, -26, -26, 71, 37, 59, -45, -3, 18, -73, 22, -37, -29, 93, -39, 13, 100, -23, -71, 29, 47, -128, 26, 124, -96, -100, 55, 70, -98, 21, 69, -90, 42, 80, -38, 38, -15, -16, 1, -127, 95, -17, 10, 5, -21, 8, -15, 1, -122, 109, 121, 37, -124, 8, 15, -128, -10, 31, 11, 74, 121, 1, -64, -85, 8, 57, -49, 34, -22, -49, -22, 58, -10, -10, 127, -22, -64, -96, -17, 93, -33, -102, 117, -24, -18, 59, -90, -26, 7, 36, 3, 11, 2, 18, -8, 53, -2, -117, 127, -23, -54, 32, -7, 37, -8, -24, -21, 64, -49, -86, 123, 102, -119, -22, 117, -53, -45, -24, -43, 97, 8, -3, -31, -29, 29, -10, 64, -29, -26, 38, 58, -70, -39, 55, -64, 43, -36, -103, 50, 44, 58, 66, 6, -65, -127, 74, 78, -128, 88, 26, -57, 80, 31, -128, -17, 15, -3, 101, 39, -86, -128, 26, 47, -26, 66, 22, -42, -11, -1, 87, 12, -48, 23, -80, 37, 102, -10, -44, -28, -15, -23, 73, 50, -6, -128, 80, 43, -58, 34, -127, 80, 73, -54, -54, -45, 127, 23, 23, -73, -90, 42, 39, -36, -93, 29, 0, 15, 127, 33, -59, -24, -66, 43, 121, -7, -65, -6, -75, -48, 127, 91, -128, -57, 127, -98, -81, 96, 81, 0, -54, -60, -63, 116, 10, -113, -5, 28, 27, 23, 60, -47, -101, 95, 108, -5, 2, -107, -59, -8, 85, 68, -15, 50, -122, -70, -15, 21, 101, 44, 17, 3, -102, -26, 70, -53, -47, 70, 97, -15, -101, 48, 28, -78, -48, 45, -26, -17, 22, 5, 103, -8, 26, -38, -128, 100, 127, -80, -36, -60, 42, 11, 27, 60, -54, -34, 43, -55, -45, 64, -76, -11, 21, 15, -7, 11, -3, -21, 33, 15, -29, -23, 15, 22, 88, -34, -90, 100, -13, -85, 13, -11, -21, 49, 127, -31, -118, -23, 45, 59, 60, -16, -97, -13, 22, 45, 59, 24, -103, -49, 33, -17, 39, 34, -78, 0, -7, -8, 59, 17, 44, 44, -12, -58, -87, -6, 93, 88, -118, -128, 54, 95, 68, 6, -113, -64, 50, -27, -6, 10, -6, -53, 127, 8, -128, 127, 3, -128, 66, -28, 68, 75, -29, -36, -11, 63, -33, 11, -34, 3, -42, 58, 0, -43, 118, -128, -34, 0, 70, 55, -69, 18, -24, 3, 34, 1, 36, -90, -15, 17, 29, 117, -6, -93, -123, 85, -8, -66, 127, 65, -47, -108, -63, 10, 36, 85, 29, -98, 21, 92, -59, -43, 28, 50, 45, 33, -93, 8, 6, -112, -43, 93, 8, -90, 44, 74, 11, -87, 38, 34, 15, 31, -66, 26, -60, -107, 74, 12, 42, 3, -127, 109, 127, -119, -109, 101, 112, -117, -128, 2, 109, 42, -2, 59, -1, -2, -76, -6, -10, -85, 31, -21, 16, 124, -13, -128, -13, 127, -16, -128, 36, 112, 71, -74, -45, 88, 2, -50, -13, 23, 53, -50, -22, 66, -128, -33, 107, -55, 47, 55, -15, 57, -8, -128, -16, 108, 18, -17, 0, -69, -45, -1, 17, 96, 24, -57, 33, -48, -71, 12, -6, 34, -26, -8, 12, -42, 8, 34, 97, -17, -50, 11, -90, 66, 49, 23, 50, -128, -42, 119, -59, -42, 49, 32, -37, 15, -33, -5, 34, 28, 17, -113, 12, -22, 68, 127, -128, -5, 16, -52, 64, 39, -39, -87, 65, 74, -39, -47, 98, -54, -78, 107, -6, -26, 32, 60, -81, -107, 17, -42, 39, 121, 28, -23, -10, 27, -91, 3, 85, -87, -8, -12, -3, 31, -45, 73, 117, -15, -128, -27, 74, -15, -88, 6, 32, 57, 57, -63, 17, -71, -75, 29, 111, 74, -127, 38, 1, -45, 81, -1, -81, 49, 127, -128, -22, 106, -127, -42, 127, -1, -116, 2, 111, -91, -96, 127, 15, -128, 42, 92, -63, 8, 22, -117, 22, 100, -15, -16, -23, -39, 45, -2, 37, 22, -18, -17, -68, 88, 43, -37, 66, -69, -45, 57, -97, -1, 127, -48, -118, 64, -18, -90, 18, 127, 7, -23, -26, -49, 111, -34, -101, -2, 44, -22, 60, -2, -103, 114, 13, -97, 16, -26, -39, 127, 26, -128, 113, 59, -92, 23, -27, -75, 127, -18, -55, 12, -95, 22, 127, 75, -31, -31, 5, 27, -65, -91, 111, 58, -96, -8, 69, -23, -24, 64, -64, -47, 111, -11, -128, 80, 69, -43, -37, 6, -24, -37, 79, 113, -98, -60, 55, -16, 11, -64, 101, 127, -90, -34, 26, -50, 55, 7, -124, -52, 90, 91, -80, -74, 90, 96, -43, -37, -18, 59, -49, -128, 127, 85, -128, 37, 55, -55, -75, 55, 12, -1, 52, -128, -11, 45, 78, -39, 36, 37, -128, 108, 127, -100, -93, 97, -53, -24, 23, -128, 121, 68, -128, 63, 127, -70, -37, -64, 59, 88, -123, -44, -37, 127, 29, -69, 38, 54, 29, -122, -79, 127, -26, -36, 95, -53, -28, -49, 38, 65, 21, -85, 7, 12, 27, 38, -48, 69, 38, -32, -118, -71, 127, 57, -128, -12, 95, 32, 52, -87, -96, 81, -34, -71, 117, 21, -128, 103, 109, -91, 33, -48, -66, 10, 81, 95, -102, -63, 2, 86, 101, -128, -33, 24, 34, 36, -78, 78, 34, -121, 31, 36, 1, -17, -68, 36, 32, -57, 3, 103, -65, 10, 21, -59, -50, -54, 45, -18, 47, 88, -97, -7, 87, 21, -65, -16, 85, 36, 12, -101, -117, 111, -6, -52, 59, 47, -16, -90, 36, 57, -3, 0, 2, -53, -8, -34, 26, 101, -111, -39, 91, 49, -42, 2, -3, -71, -8, 49, 98, -79, -43, 108, 58, -123, -8, 24, 18, 44, -7, -17, -2, -50, -17, 80, -47, 29, -11, -122, 59, 127, 8, -91, -2, 12, -8, 2, -39, 0, -76, 86, -11, 23, -3, -80, 127, 71, -47, -58, -75, 12, 22, -57, 10, 5, -10, 102, 27, -128, 73, 27, -18, 102, -52, -85, 73, -36, 6, 111, -15, -93, -21, 18, -33, 69, 44, 15, -57, -6, 7, -73, 0, -55, 87, 65, -80, -70, 63, 81, -127, -3, 127, 43, -128, -2, -11, 48, 64, -123, -34, 97, 116, -64, 5, 55, -113, -52, 127, -39, 1, -1, -74, 112, -90, -101, 95, 97, -74, -33, 78, -22, 3, 38, -80, -107, 34, 114, 88, -106, -90, -8, -16, 107, 1, -21, 6, 26, 58, -42, 33, -11, -49, -12, -22, -27, 53, -28, 1, 121, -45, -11, 91, -103, -33, 53, 6, -34, -33, -17, 0, 127, -5, -15, -95, -29, 119, -7, 23, 0, -54, -24, -28, 27, 17, 10, -50, 2, 85, 16, -13, -42, -86, -42, 8, 76, 127, -48, 6, 71, -116, 28, 93, -128, -96, 127, 98, -26, -128, -23, 75, 10, -74, 3, 24, 0, 113, 21, -60, -106, -63, 66, 1, 54, 87, -12, -21, -65, 23, -36, -70, 28, 13, 95, -18, -45, 16, 36, -54, -85, 66, -34, -65, 91, 86, -43, -80, -12, 127, -73, -49, 127, 42, -102, -8, -28, -97, 60, 80, -57, -107, 101, 65, -92, -31, 32, 48, -10, -59, 42, -29, 37, 127, -6, -128, 11, -24, 15, 109, -66, -96, 44, 95, -71, -3, -48, 36, 10, -111, 127, -23, -42, 127, -1, -119, -86, 95, 36, -118, 24, 73, -15, -7, -10, 69, 55, -128, 21, 63, -128, 100, 53, -107, -57, 58, 44, -32, 47, 71, -66, -123, 79, 107, -13, -57, -74, 33, 53, -8, -21, 52, -17, -128, 81, 127, 22, -93, -73, 18, -44, 6, -33, 80, 96, -127, 68, -47, -53, 74, -1, 50, -93, 3, 17, -91, 118, 47, -23, 17, -48, -79, 58, 93, 0, -18, 0, -26, -118, -53, 85, -15, 37, 100, -127, 71, 23, 10, -27, -116, 69, 45, -15, -24, 42, -78, 43, 100, -128, 54, 8, -128, 18, 127, -58, 31, 36, -128, 127, 33, -11, -39, -70, 91, 42, -64, -93, -2, 127, -39, -90, 93, 45, 15, -26, 3, -90, -85, 114, 34, -80, 29, 55, -92, 23, 70, -31, 49, -80, -59, 76, -18, 48, 97, -22, -16, -97, -38, 74, -81, 10, -1, 12, 127, -54, -66, -15, -68, 27, 15, 63, 86, -18, -80, -65, 121, 39, -108, -8, -48, 48, 59, -78, -70, 122, 127, -128, -47, 101, -12, 8, 36, -11, -55, -28, 43, -60, -10, 86, 1, -85, 32, 10, -92, 96, 74, -2, 39, -128, -11, 98, -78, -33, -53, 66, -1, -29, 64, -68, 92, 26, -128, 38, 111, -39, -55, 49, -24, 33, 103, 0, -60, -39, 18, 54, -54, -45, 43, -42, -55, 80, 12, -118, 85, 127, -65, -87, 43, -55, 10, 127, -15, -128, -53, 122, 95, -57, -18, -26, -116, 59, 127, -98, -96, 54, 81, -16, 6, 21, -118, 8, -18, -11, 102, -27, -121, 87, 23, -57, 90, -8, 29, -42, -76, 76, 70, -57, 11, 27, -98, 15, 118, -60, -111, 1, 29, 2, 22, 119, -21, -53, -32, -79, 36, 113, 18, -95, -7, -2, -12, -1, 55, 16, -81, 92, 37, 10, -39, -45, -39, -78, 85, 73, -3, -64, -74, 127, 8, -29, 29, 27, -11, -97, -31, -29, 127, 23, -52, -12, -57, -31, 58, 127, -43, -91, 80, -87, 18, 109, -112, 50, 42, -24, -38, -1, 8, 34, -32, 3, 81, -10, -88, -71, 23, 95, 15, -106, 3, 63, 76, -85, -6, 79, -38, -79, -29, 113, -22, 3, 55, -45, -69, -96, 118, 76, -108, 65, 16, -48, 65, -16, 8, 54, -48, -81, 68, -10, -78, 75, -34, 7, 113, -106, -111, 63, 36, 53, 71, -88, -69, 69, 34, -53, 36, 45, -60, -23, 52, 22, -128, -101, 22, 127, -39, -53, 127, 3, -92, -7, -49, 47, 76, -128, 97, 68, -44, 60, -88, -79, 90, -16, -64, 5, 38, 44, -57, 69, -37, 6, 66, -69, -8, -80, 78, 85, -71, -21, -29, 53, 53, 5, -47, 1, 63, -65, 55, -48, -90, 127, 0, -119, 50, 38, 5, -11, -24, 18, -87, -37, 60, -24, 43, 26, -15, 29, 3, 18, -38, 59, -55, -122, 18, 50, 15, 12, 63, 50, -121, -87, 100, -26, -12, 111, -88, -60, 127, -24, -34, -3, 32, 2, -85, 5, 97, -39, -64, 45, 31, -42, -74, 3, 111, 38, -124, 17, 2, -26, 79, -45, 3, -8, -76, 127, 42, -128, -10, 68, -37, 11, 29, -53, 55, -31, -23, 91, 24, -81, -80, 79, 54, 75, -88, -74, 98, 37, -24, -111, 16, -6, -1, 127, -73, -34, 52, 8, -42, 18, 112, -13, -128, -71, 15, 39, 53, -12, -50, -29, 55, 39, -79, 66, 95, -23, -68, -68, -24, 108, 12, -127, -8, 69, 127, -2, -95, -47, -49, -18, 127, -39, -10, 22, 2, 92, -33, -27, -6, -36, -76, 59, 60, -100, 7, 127, 33, -32, -8, -36, 37, 27, -43, -90, -23, 16, 29, 114, -6, -128, 10, 96, 23, -70, -90, -31, 106, -11, -60, 127, 38, -55, -73, -60, 76, 48);
 
    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project
 
    constant SCENARIO_ADDRESS : integer := 100;
 
 
    --Scenario 2
    constant SCENARIO_LENGTH2 : integer := 12000;
    constant SCENARIO_LENGTH_STL2 : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH2, 16));
    type scenario_type2 is array (0 to SCENARIO_LENGTH2-1) of integer;
    signal scenario_config2 : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
    to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
    1,                                               -- S
    0, -1, 8, 0, -8, 1, 0, 1, -9, 45, 0, -45, 9, -1           -- C1-C14
    );
    signal scenario_input2 : scenario_type2 := (50, 99, 107, 1, -120, 36, 3, 28, 6, -109, 81, -109, 60, -29, 65, 65, -107, -117, -19, 48, -95, -38, 86, 80, 31, -29, 29, 1, 87, -122, -105, 42, -36, -80, 0, 79, -117, -37, -79, -109, 120, 35, 62, 70, -71, -36, 10, -65, -71, -7, 44, -47, 91, -86, -19, 118, -75, -60, -114, 26, -125, -97, -8, -124, -73, 52, 123, 88, -39, 122, -27, 0, 47, 66, -35, 91, 107, 103, -80, 127, 88, -50, 73, 126, 121, -128, 103, 92, 59, -107, -71, 74, 8, -115, -96, 13, -116, -59, -99, 93, -46, 82, 3, -83, 101, 30, 110, 41, 88, -101, -64, 115, 45, 117, 58, -25, -57, -52, 108, 118, -24, 29, -106, 3, 52, 84, -53, -82, -75, 27, -41, 15, -122, 93, 77, 106, -10, -73, 37, 20, 35, 67, 12, 51, -39, -83, 93, -79, 111, -68, -94, 6, -55, 91, -126, 67, -14, -72, -7, -62, 0, -54, -36, 108, 54, 121, 64, 37, -13, 58, 96, 36, -32, -91, 121, 102, -89, -32, 125, 114, 71, 72, 29, 89, -47, 79, -20, 20, 74, 1, 101, -127, 15, 13, -88, -107, -59, -57, -84, -1, 21, 8, -37, 118, 26, 122, 69, 6, 111, 74, 32, 73, 34, -56, -53, 82, 72, -87, 39, -119, -23, 94, 93, -95, 69, 118, -72, -45, -64, -99, 118, -39, -78, 83, 75, -27, -104, -43, 85, 124, -57, -43, 76, -32, 5, -53, 9, -72, -52, -86, -9, 54, -97, -46, -13, 21, -67, -127, 3, 86, 6, -94, -31, -10, 120, -52, 70, -68, -116, 114, -27, -113, 14, -45, -82, 116, 15, 111, -110, 76, -98, -87, 109, -67, 86, 86, 8, 13, -10, -24, -48, -110, -106, 8, 109, 30, -43, 108, -90, 38, -53, -101, -37, -15, 6, 54, 0, 108, -43, -102, -3, 116, 103, 116, 48, 86, 122, 119, -104, -6, 67, 95, -50, -115, -62, 73, -101, 4, 127, 13, -25, 71, -90, -83, -5, 122, -22, -112, -117, -11, 86, 59, 46, 10, 123, 47, -48, 11, 5, 40, -4, -6, 3, 104, 105, 39, -62, 27, -64, 65, -67, 0, -123, 86, 57, 13, -1, -27, -43, -16, -70, 63, 127, 107, -111, 59, -57, 28, 0, -81, 0, -75, -54, 28, -58, -36, -78, -94, 21, -13, -26, 3, 11, -20, 126, 127, 47, -5, -67, -101, -27, -57, -96, 56, -93, 51, 21, 105, -107, -31, -72, -66, -118, 96, -8, -47, 114, 116, 70, -15, -54, -97, -82, 115, -38, -16, 25, -67, 95, -38, -54, 89, -121, -61, -87, -9, -107, 66, -6, 77, 84, 42, -108, -27, 65, -121, 123, 36, -71, 69, 9, -51, -24, -116, 47, 108, 72, -107, 62, 120, 13, 125, -77, -80, 120, 116, -41, 66, 60, 61, 65, 0, 113, -2, 65, 24, 116, 48, 105, -3, -53, -68, 72, 67, -106, 101, -113, 74, -122, 14, 46, 115, 48, -80, -39, 80, -126, -127, -21, 58, 97, 102, -107, -12, -92, -21, 35, 9, -3, 53, -17, 13, -92, -42, -118, -32, 117, 12, 57, -122, 94, -20, 116, 39, 37, 69, -126, 83, -71, 51, 4, 81, 121, -48, -43, -5, -65, -9, 41, 112, -41, -126, 43, -2, -115, -124, 121, 101, 63, -82, -12, -88, 13, -98, 108, 110, 66, -4, -15, 74, -14, -45, -67, -67, 124, 98, 14, -92, 84, 93, -71, -123, 62, 40, 100, -52, -50, -74, 113, 42, 42, -23, -3, 45, 94, 65, 17, 64, 84, 79, 68, 99, 110, 98, 108, 73, -52, 17, -93, -61, 123, 11, -49, -76, -78, 117, -51, -126, -118, -36, -24, 92, 117, -3, 105, 98, 62, -43, 56, -67, 16, 27, -37, -128, 15, -16, 34, -40, 39, -25, 27, -74, 84, 105, 24, 25, 33, -81, 96, -36, -23, 48, 55, -49, 53, 78, -107, 110, -35, -97, -63, -35, 65, 42, -118, -96, 12, 48, 114, 76, -44, 30, -22, 53, -73, 14, -33, -97, 50, 31, -1, -30, -25, -11, 0, 104, -102, 111, 95, -1, -78, 24, -109, 60, -22, 11, 23, 71, -42, -2, -84, -73, 90, 74, 21, 31, -84, -84, 24, 105, -6, -58, 31, -80, 15, 124, -109, 15, 83, -18, 109, 64, 17, 45, 109, -8, 108, 85, 108, 84, -90, -41, -83, 78, -19, -110, 23, 61, -19, 110, 36, 63, -13, 18, -105, 3, -91, 9, 59, 8, 6, 110, -114, -39, -31, -71, -10, 34, -37, -11, -6, 83, -10, 107, 113, 52, -3, 15, 27, 0, 74, 45, -89, 34, -106, -102, -66, 51, -63, 76, -126, -19, -47, -17, -112, -29, -109, 35, -9, -59, -25, -97, -104, -54, 2, 107, -89, -81, -115, 111, 127, 55, -5, -97, 100, -81, -125, 109, 48, -41, -118, 41, -128, -126, 71, 37, 3, -45, 5, 94, 65, 63, 95, 19, -42, 82, 23, 97, 75, 54, -14, -25, 117, -38, 83, 77, 97, -95, -71, -26, -120, 108, 3, -78, 115, 33, -7, -20, 13, 94, -102, 65, -42, 126, 115, -81, 2, 36, -20, -103, -41, 77, 12, 121, 33, 111, 20, 6, 6, -124, -77, -44, 117, -24, -22, 94, 10, -109, 12, 5, -43, 0, -120, 61, -110, 105, -87, 22, 5, -54, 94, 78, -108, -122, -11, 51, 45, 51, 45, 113, -14, 12, -7, -109, -5, -90, -81, -121, 13, -44, -65, -65, 60, -110, -89, -20, 57, -4, -21, -24, -54, -65, -126, 110, -39, 14, 43, 20, 19, 10, 64, -45, 50, 109, 35, -101, 106, -83, -94, -110, -64, -68, -6, 88, -96, 48, 93, 21, -88, -42, -1, -64, 41, -127, 7, -24, 58, 7, -38, -34, 27, 42, 59, -50, -2, 69, -124, -29, 20, -55, 23, 41, 82, -21, 53, -51, -48, 125, -39, 19, 41, 98, -111, 8, -117, -96, 74, 41, 60, -65, 38, 31, 3, -18, 26, -68, 108, 85, -56, -2, 42, 100, -113, 114, 85, -16, -55, 77, -65, 46, -107, 76, -37, 36, -10, -22, 44, -39, -88, 73, -120, -42, 89, -20, 102, -96, -65, 53, -58, 106, 47, -60, 100, -27, -15, -15, 16, -98, 38, -64, -47, -12, 111, 17, -46, 91, -44, -68, 21, 4, -115, -108, -55, -62, 103, 78, 18, -115, -108, 105, -19, -14, 81, -125, 115, -123, -108, -28, -20, -125, -32, 62, 77, -44, 14, -46, -61, -8, -52, -10, -42, 54, -86, 49, -18, 97, -77, -113, -4, 105, -77, -112, -125, -15, -8, 48, 23, -84, 2, 22, 112, -32, 118, -24, -73, 28, 69, -126, 86, -115, -76, -104, 111, 36, 60, 59, 41, -33, -83, 45, 56, -100, -31, 119, 92, 112, -18, -78, -35, -113, 2, -128, 88, -23, 122, 110, 26, -57, 35, 29, -95, 48, -51, 101, -113, -23, -46, 109, -118, -86, 64, 32, 61, 90, 126, -37, 48, -21, -13, 107, -107, 37, -5, 56, 91, 18, 87, -72, 85, 36, 76, 81, 25, 40, -114, 62, 19, 39, 24, -26, -112, -5, -73, 10, 75, 31, 108, -52, 50, 44, 69, -18, 113, -128, -11, -98, -15, 49, 85, -103, 84, -60, 30, -61, 40, 77, 40, 76, -81, 93, -17, 67, -48, -30, -107, -8, 104, -77, -85, -10, -37, 24, 69, 123, 85, 74, 34, -85, -113, 79, 123, -111, 51, 55, -34, -99, 117, -14, -4, 70, 13, -39, -41, -60, -40, -99, 76, -49, -9, -110, 53, 118, 2, 65, -88, -77, -13, 126, -121, 120, 66, 67, 19, 93, -114, 99, -120, -84, -96, 99, 72, -101, -20, 94, 24, -111, -36, 4, 55, -96, 121, -108, -60, -121, 43, -106, -96, 103, -97, -127, -14, 94, 102, -6, 79, 91, -30, -45, -127, 84, -68, -57, -88, 125, -127, 59, 34, 39, 87, 71, -30, -32, 66, -102, 79, -51, -126, 2, -5, -123, 47, 71, -105, 21, -103, 67, 97, -71, 22, -107, 96, -44, 30, -21, 47, -35, -127, -89, -109, -11, -56, 120, -118, -115, -53, -21, -8, 112, 88, 71, 110, 124, 75, 77, -92, -35, 86, -11, 47, 94, 121, 94, -39, 47, 121, 127, -45, -46, -66, 60, 51, 109, 17, 108, 88, 51, 33, 57, -114, 15, 36, -6, -38, -91, 20, -37, -95, -6, -27, -19, 15, -78, 77, 107, 112, 47, 122, 70, -11, 64, -71, -11, -72, -13, 25, 120, 118, -13, 29, -113, 21, 18, -73, -59, -34, -5, -24, 22, -110, 123, -128, -81, 81, -45, -35, 67, 0, 86, 55, -16, 0, 109, -119, 100, 62, 16, 75, -47, 84, 15, 37, -103, 81, -9, -125, 98, 39, 86, -102, -36, 122, -74, -6, 93, -112, -80, 47, -55, -28, -42, -126, 80, -63, -34, -13, -80, 51, 105, 43, 34, 20, 36, 0, 47, 123, -106, -117, -81, 118, -60, -54, -30, 34, 13, 8, 107, -62, -41, 29, -39, 48, -126, 46, -111, -3, 114, -9, -23, 125, -88, -73, 122, -48, 93, 37, 72, -32, -16, -59, 67, 63, -120, 10, -22, -81, 95, 120, -46, 102, -79, -93, 79, -43, 100, 4, 108, -112, 86, 117, 35, 36, 123, 125, 2, 116, 76, 108, -50, -82, 47, -18, -23, 92, -11, 101, 21, -93, 50, -36, 71, 32, -54, -74, -88, 76, -109, 78, 69, 41, -80, 1, 4, 61, -19, -72, -13, 111, 102, 46, 91, 93, -92, 15, 6, -120, -19, 68, -111, -45, -58, 88, -21, -30, -56, 79, 84, 44, 87, -108, 80, 88, -85, -84, 72, 87, -85, -19, -128, 100, -104, -126, -28, 85, 124, -28, -59, -10, -51, 19, 0, -100, -34, -1, -107, 28, 56, 97, -46, -43, 109, 59, 120, -114, 102, 53, -42, 42, -36, 27, -30, 79, 60, -60, 90, -8, -88, 52, -66, 62, 116, -76, -53, 75, -40, 16, 19, -21, -65, -62, 86, -38, -66, -31, -20, -72, 62, -26, 42, 110, -57, 50, -62, -110, -43, -73, 101, -44, 80, 29, 83, -94, -36, -73, -122, 112, -73, 13, -102, 115, 37, 27, -85, -96, 126, -6, 109, -67, -122, -20, -43, 102, -17, -95, -60, -120, -14, 77, -6, 120, 79, 13, -120, -121, -27, 110, -23, -92, -20, -124, -99, 20, 78, -99, -121, -51, 23, -49, 109, 91, 87, 67, 4, 82, 26, -107, 27, 65, 19, 18, 60, 50, -37, 64, 91, 35, -3, -113, 55, -93, 120, -4, 79, 105, -29, 99, 71, 64, 83, 84, 21, -35, -29, -107, 35, 95, -38, 73, 76, -105, 79, -112, 8, -116, 95, -50, 24, -55, -72, -76, 43, -8, 118, 87, 84, 95, -59, -4, -20, 115, -66, -90, -105, -95, -47, -89, 106, 66, -81, 100, -42, 68, 110, 126, -88, -1, -90, -92, 33, 72, 74, -102, 87, 102, 26, 19, -56, 121, 8, 63, -87, 127, 34, 14, 86, 112, 91, -51, -34, 24, 112, -39, -32, -50, -101, 9, 65, 73, 18, -20, -80, -85, 87, -34, 73, -3, 109, 79, 122, 92, -42, -115, 37, 26, -115, 23, -38, 68, 75, 90, 82, 108, -39, -94, -36, -62, -36, 1, 52, -38, -123, 83, -75, -59, -48, -13, 88, -56, 66, -112, 76, -14, 58, 61, -86, -15, -43, 12, 25, -111, 124, 46, 5, -47, 115, -90, 97, -101, 50, -40, -116, 86, -127, -101, 49, 48, -37, -28, -35, 13, -91, -7, -16, -42, -83, -66, -81, -36, 10, -110, -124, -77, 34, -98, 1, -55, 108, -20, 27, 67, -62, -61, -53, -87, 110, 22, -81, -56, 17, -86, 16, 34, 68, -49, 126, 51, 41, 85, 124, 116, -122, -109, -60, -79, 54, 126, 30, -16, -86, 14, -91, -83, -43, 53, -120, -13, -72, -49, -53, -11, 56, 62, 92, 43, 35, 68, -35, 114, -52, 8, -22, -3, -92, 102, -77, 36, 92, -21, 87, 49, 59, -112, 0, 20, -25, -106, 18, 46, 69, 50, -80, -71, 49, -7, -3, -47, 64, -72, -104, 121, -14, 37, -98, 95, 115, -111, -47, 82, -114, -38, 84, -29, 107, -77, 73, -20, 92, -13, -3, 123, 0, 64, 22, 0, 73, -43, -65, 103, 51, -117, -29, 28, -7, 75, 28, 90, -54, 66, -109, 102, -28, 45, 8, 31, -90, 47, -87, -2, -91, 115, -90, 67, -39, -119, 23, 113, -23, 14, 5, 56, 77, 51, 108, 93, 52, 97, 120, -63, -79, -66, 91, 124, 106, -35, 16, 28, -106, -124, -18, 35, 47, -46, -117, 109, -37, 5, -49, 4, 38, -97, 38, -57, -105, -16, -118, 105, -103, 37, -29, -40, -16, -70, -28, 53, -111, 26, -83, -116, -128, 46, 32, -49, -124, 100, 33, 48, -75, 74, 17, 24, 56, -24, -100, -61, -19, 9, 101, -22, -90, 85, -9, 2, 120, -83, 36, -82, 91, -114, 73, -40, 115, 39, -13, 34, -101, 47, 74, -51, 57, 125, 123, 85, -74, 14, -1, -62, -66, 89, 89, 79, -69, -90, -85, 80, 37, 83, 72, 48, -68, 22, -115, 1, -71, 10, -108, 38, 42, 12, -125, -122, -8, -82, 67, -51, -47, -1, -80, 90, -42, -91, 97, -63, 18, 61, 15, 125, -83, -13, -16, 8, -52, -88, 1, -57, -127, -33, 48, -47, -120, 106, 106, 120, 31, -89, -3, -52, 36, 14, -109, 52, -107, 89, 62, 105, -20, -38, -64, -77, 110, -123, -89, -22, 79, -115, -9, -37, -112, -126, -71, -87, -79, 64, -3, 43, 33, -26, 122, 114, -76, -40, 8, 11, -73, 62, -119, -95, -15, 28, 119, -38, -39, -75, 26, 57, -69, -78, -93, -43, 94, -96, -59, 83, 99, 57, 124, -8, -51, -18, 22, -113, -41, -27, -79, 16, 5, 26, 96, -114, -70, 49, 107, 84, -58, -109, -53, -104, -11, -70, 97, 65, -11, 104, 54, -34, 85, 18, 124, 47, -18, -4, -97, -124, -111, -94, 126, -103, 109, -53, -67, -102, -46, -127, -122, 79, 19, -103, 58, 120, 13, 103, -55, 19, 122, -64, 103, 27, -118, -1, -6, -5, 69, 113, -22, -124, -29, 72, 73, -45, -37, -29, -117, -80, 57, -6, -41, 74, 69, 112, -82, 31, 38, -96, -121, -119, -116, 16, -10, 93, 73, -71, -93, -23, 114, -1, -35, -103, 69, 123, 0, -122, 112, 28, 109, 120, 57, -45, 50, 98, -47, 37, 104, 7, -97, 107, 23, -74, 65, 31, 121, 78, 15, 58, -64, -103, -1, 97, -100, 123, 27, 58, -94, -103, 13, 30, -116, -17, -99, -87, 39, -44, 98, 120, -53, -65, 38, -37, 88, -107, -23, -22, 25, -31, -87, 125, 54, 91, -111, 69, 32, -95, 24, -100, 30, 92, -101, -40, -39, -93, 47, -100, -71, -22, 68, 66, -89, -36, -89, 69, -127, 58, 95, -31, 125, -31, -55, 50, -119, 74, 25, -128, 89, 21, -106, -122, 79, -61, 123, -116, -4, 64, 38, 55, -116, -76, 31, -58, 41, -40, 26, -79, 48, 59, -49, -98, -4, 95, -55, 26, -35, 11, 33, 8, 10, 110, 109, -100, -36, -95, 63, -81, 69, 108, 74, -2, 74, 67, 89, -79, -101, 30, -37, 57, -20, 101, -66, 57, -15, -42, 49, -36, -7, 76, -16, 76, -17, -15, 67, 47, 37, 115, -26, 114, -90, 83, -37, 74, -109, -100, 33, 18, -12, 119, 73, 88, -114, -107, -25, 102, -36, -27, -13, 97, -82, 115, -7, -76, -78, 121, -23, -11, -41, -35, 116, -105, -61, 93, 44, 50, 116, -95, -97, 85, 113, -118, 80, -127, -63, 117, 116, -8, 80, 23, 1, -40, 45, 70, 27, -73, 91, -110, 0, -106, 53, -110, 123, -30, -9, -33, 9, 8, 104, -57, -121, 103, -64, 14, 82, -80, -50, -25, 46, -41, -20, -14, -16, 98, -26, -123, -32, 76, 101, 16, 54, 100, -35, 114, -36, 46, -30, -82, 45, 94, -124, -30, -27, -86, -38, 83, 10, -117, 25, -44, 4, -109, 51, 104, 81, 99, -91, 64, -60, -5, 59, -43, -21, -25, -5, 33, -27, -65, -66, 110, -102, 70, -87, -110, -74, 28, -16, 74, 116, -71, -95, -61, 96, 56, 44, 85, -55, 124, 55, 63, -56, -95, -81, -83, -73, 75, 123, 71, -110, 74, -64, -76, 24, -7, -122, 112, 65, -112, -30, -74, 58, 30, 111, 76, 81, -124, 16, -30, 5, 119, -60, -3, -38, 11, 107, 72, -99, 124, 29, -28, -55, -62, -98, 87, -122, -19, -81, 95, -107, -19, 94, 125, -101, 87, 65, -110, 4, -5, -21, 69, 48, 22, 58, -9, 85, -114, -91, -29, -123, 22, 36, -45, -112, 66, 13, -50, -83, -111, -62, -58, 41, -118, -67, -84, -126, 88, -127, -42, 5, 82, -15, 71, 27, 43, -31, 106, -93, 10, -109, 12, -15, -19, -119, 33, -106, -122, 53, -78, -47, 31, 17, -105, 53, 120, -109, 80, -110, -55, -55, 79, 124, 45, 6, 66, -60, 39, -44, -27, 26, -87, -106, -55, -96, 50, 59, -58, -128, -7, 36, 90, -66, -39, -35, -94, -89, 69, -123, 66, 125, -102, -98, -63, 100, -90, -102, 61, -113, 113, -65, 109, 90, -115, -99, -83, -101, 44, 2, -83, 97, 42, -120, -54, -91, 96, -7, -17, -23, 122, -36, 15, 96, 48, 125, 40, -87, 63, -71, 110, 4, -80, 40, 25, 125, -19, 5, -23, -2, -13, -34, -123, -74, 12, -13, 27, -22, 80, 7, 122, -83, -10, -124, 62, 21, -22, -21, -104, 47, -46, 120, -55, -32, -32, -14, 119, 118, 81, 77, 78, 106, -16, -36, 37, -69, 127, -15, 46, -31, -73, -1, 34, 53, -43, 7, 33, 111, 77, 96, -102, -46, -62, -4, -83, 22, 55, -85, 122, 110, 89, 103, -7, 103, 120, -25, 46, -126, 69, -31, -4, -65, 126, -24, -5, 126, -71, 79, -94, 49, -53, -104, 99, 23, 35, 82, 8, -6, -102, -16, 74, -49, 51, -88, 9, -16, 46, -87, 43, -45, -73, 103, -111, -79, 101, 55, 80, -89, -74, -85, 121, 36, 96, 97, 50, 7, -32, 70, -87, -127, 49, 6, 41, 83, 78, 62, -54, -106, 34, -41, 59, -45, -115, -3, 35, -15, -87, 79, 83, 90, 14, -13, 71, 25, 87, -42, 19, 70, 60, 72, -93, -25, -106, -82, -96, -36, 30, -104, -36, 84, 37, 122, -125, 123, 61, -79, -99, -87, -36, -65, 105, -83, 38, 54, -84, 52, -94, -71, -100, -32, 91, 7, 8, -87, -46, 111, 59, 97, 84, 92, 88, -76, -93, -25, 25, -128, 26, 57, 21, -16, -54, -126, 35, 111, -45, 17, -9, 54, -31, 73, 42, 74, 2, 7, -13, 99, 4, -61, -32, -23, -101, -60, -21, 25, 60, 26, -58, -105, 0, 62, -8, 70, 17, -91, -52, 62, 104, 17, -16, 85, 4, -122, 16, 99, 3, -60, 108, -102, 64, -53, 123, -91, -99, -32, -98, 122, -74, 81, -36, -36, -102, 9, 82, -105, 45, -24, -104, 109, 119, 78, 124, 64, 14, -16, 90, -34, 39, -80, -24, 114, -44, -27, 29, 125, 95, -52, 34, 86, -10, 82, 53, -115, -128, 20, -124, -65, -46, 77, 62, -50, -108, -22, -77, 121, -72, 36, -65, -15, -98, 119, -92, 84, 12, 10, 10, 78, 98, -124, 31, -79, 71, 43, 10, -64, 91, 105, 61, -55, -94, 63, -46, -93, -77, -20, 27, 48, 106, -19, 99, -94, -71, 87, -96, 124, 43, -23, -126, 7, -75, -31, 67, -10, 83, -12, -62, 92, -50, 38, 72, 60, 68, 43, 93, 24, -2, 96, 7, -30, 106, 47, -40, -120, 84, -113, -23, -21, -78, -106, -89, -53, 36, 50, -13, 50, 47, 13, -36, 65, -62, 71, -54, -85, 54, -118, -128, -63, 84, 33, -49, -87, -41, -85, 50, -35, -70, 106, 76, 1, 26, 94, 54, 59, 63, -67, 92, 78, 87, 92, -16, -112, -35, 108, -94, 21, 97, -114, -51, -62, -88, 53, -64, -80, 36, 18, 31, 57, -90, 120, 20, 115, 52, 6, -44, 64, -71, -34, 49, -67, 78, -43, 99, -126, 77, -60, -2, -2, 44, 113, 83, -7, -28, 67, 102, -124, 54, 29, -105, 84, 8, 120, -11, 12, -85, 100, -43, 38, 37, 48, 15, 88, -48, 66, 98, 62, 15, 91, 109, -83, -75, -15, -16, 75, 65, -3, 43, 41, 73, 102, -94, -115, 81, -110, 127, -71, 87, 79, -40, -19, 61, -112, 64, 50, 88, 28, -47, -123, -125, -78, 79, 39, -24, -6, 59, -62, -92, -4, 114, -57, 21, 3, 39, -82, -76, -112, -8, -21, 90, -74, -52, -86, 102, -103, 123, -105, 61, 124, -62, 97, -69, -101, 50, 9, 57, 121, 23, -57, 56, -66, -69, -9, 29, -92, -12, -69, 23, 67, 16, -77, 125, -46, -44, -55, 25, -56, 108, -108, -98, 43, -64, -77, 47, -124, -123, 59, 49, 84, -70, -31, 125, 61, -14, -6, -110, 98, 57, -10, 59, 87, -77, -37, -128, 102, -22, -128, -9, 59, -18, 96, 79, -95, 87, 35, -11, 87, -45, 94, 20, 14, 117, 93, 28, -54, -28, 102, 81, 52, 98, 83, -104, 36, -109, 47, 119, -119, 101, 64, 101, 109, 72, 19, 80, 121, 22, -2, -74, 81, 121, -74, 47, -64, -73, -63, 50, -93, 40, 7, 50, 108, 124, 39, 125, -77, 21, -85, -63, -25, 47, 104, 18, 42, -124, -46, 66, 51, 112, 20, -15, -31, 70, -102, -34, -45, -62, -116, 33, -117, 42, 89, -20, -24, -79, -45, -35, -15, -90, 72, 76, -72, 99, -17, -44, 2, -115, 80, 77, -6, -24, -8, 53, 119, -111, -36, 44, 99, -86, 44, -108, 31, -18, 48, -96, 104, -55, -6, -42, -72, -112, -9, -118, 28, -37, 46, 73, 67, -79, -72, -116, 33, 75, -100, 125, 84, 114, 10, 100, 109, 52, 27, 70, 48, -82, -36, -22, -57, 127, -84, -32, 57, 118, 71, -2, 2, -112, -121, -60, 32, 40, 82, 23, -32, 44, 70, 13, 111, -85, -42, 3, 12, -7, 33, 37, 21, 58, 61, -41, -55, -105, -34, 49, 42, -75, -14, 109, 114, -93, -89, 105, 91, 58, 72, 95, 122, 13, 53, 110, -4, 36, 62, -111, -79, -79, -95, -67, -55, 125, 67, 104, 10, 9, -126, -26, -127, -105, 24, 96, -108, 85, 38, 84, 3, 65, 112, 24, -72, 67, -3, -72, -75, -66, -99, -32, 61, -49, -79, 8, -114, -15, 5, 69, 119, 55, 118, -97, 84, 126, 122, -97, 62, 22, -22, -65, -40, 0, 35, -74, -114, -127, -72, -96, -104, 41, -35, -23, -2, 95, -77, 83, 12, -7, -4, 126, -95, -57, 121, -77, 17, 26, 114, 84, 102, 91, -68, 93, -108, 103, 6, -60, -83, 111, -88, 37, -48, -108, -114, -88, -59, 40, 72, 97, 42, 116, -78, 2, 120, -32, -5, 65, 8, -108, -74, 76, -17, 117, -2, -78, 22, -37, -90, 60, -111, -106, 4, 119, 78, -40, 51, 77, 56, 89, 51, 12, 0, 117, -29, 38, -32, 73, -76, -61, -76, 106, -109, -119, -57, -104, 52, 51, -121, -36, -117, 80, 28, 71, -105, -127, 126, 23, 61, 111, -63, 4, -73, 86, -79, -81, -117, 102, -108, -91, -52, 7, -60, -38, -124, 91, 76, -3, -19, 27, -100, 2, -105, 2, -97, -7, -80, 100, 19, -35, 87, -23, -19, -79, -63, -15, -37, 22, -111, -65, -75, -98, -96, -85, 80, 13, -40, -70, 115, -109, 89, -93, 111, 8, 1, 21, 50, 108, -52, -123, -66, 5, 28, -26, -7, -11, -107, -49, 86, -103, 81, -28, 41, -24, -15, 112, -53, -91, 13, -28, 45, -80, 5, 107, -51, 31, -82, -114, 24, -123, -27, 106, 127, -27, 93, -11, -34, 47, -108, -118, -125, -19, -72, -61, 53, -31, -87, -82, 70, 122, 20, 78, 29, -1, 52, -67, 9, 25, 16, -26, -14, 94, -123, 36, 56, -70, -29, -104, -8, 24, 11, -17, 80, -79, 14, -25, 31, -118, 55, -96, -106, 1, 34, 36, 101, 115, 56, -27, -28, 2, 99, -102, -34, -86, -79, -28, 86, 17, -89, -85, 11, 8, -115, 1, -108, 80, 38, -106, -60, 114, -70, 85, 111, 47, -59, -124, -48, 103, 76, 46, 5, 95, -41, -122, -39, -72, -102, -99, 2, 70, 27, 112, 32, 7, 106, 4, 114, -107, 86, -45, -38, -8, -100, 29, 100, -128, 66, -112, -71, -47, 18, 63, 127, 4, 10, 23, -32, 107, -5, 78, -25, -53, 36, 101, 20, -68, -95, -26, 43, -21, -39, 86, -26, -119, -8, -9, -9, 90, 17, 103, 26, -84, -59, -33, 89, -27, 19, 38, 86, 27, 77, 27, -22, -22, 10, -96, -112, 77, -63, -37, 17, 123, 36, -113, 26, -122, 60, 122, 45, 91, -106, 13, -104, 84, -66, -48, -98, -10, -13, -127, 25, 0, -17, -91, 19, -80, -114, 64, -102, 29, 7, -20, -31, 47, -112, -11, -59, -97, 88, 46, -4, -52, 9, -4, -120, 75, 61, -97, -121, 63, -18, -20, 52, 45, -96, -64, 63, 45, -8, 118, 75, -107, 70, 79, 21, 72, 69, -94, 81, 63, -101, 10, 124, 20, -104, 16, -98, 58, 100, 120, 33, 44, -103, -72, -112, -53, 44, -110, 76, 1, 79, 71, 44, -22, 114, -123, -12, -110, -50, 106, -20, -111, -24, -116, 58, -60, -27, -31, -94, -10, 45, 120, 6, 71, -15, -120, -17, -89, -12, -75, -29, 119, 34, 70, 100, 57, 60, -94, -57, 95, 113, -29, -40, -94, -75, -115, -91, 17, 60, 121, -48, -37, 20, -37, -8, -90, 69, -21, -91, 84, -33, -98, -26, 98, 75, 29, -34, -37, -73, 69, 54, -18, -12, 3, 115, 76, -50, -125, 77, -8, 18, 31, 40, 15, -109, -9, -24, -126, 19, 32, 124, 56, 43, 2, -97, -92, -87, -17, 65, 70, 94, -106, -115, 19, 7, 113, -53, 37, 20, 117, 0, -75, -64, 111, -20, -78, -13, 82, 109, -105, 82, -89, 55, -101, -29, 65, -91, 44, -92, -23, 54, 31, -37, 75, -107, -41, 18, 101, 117, 120, 17, 89, 32, 58, 114, 48, 33, 74, -126, -70, -92, -30, -72, 107, 44, 119, -37, 124, 118, -36, -1, -14, -84, 96, -4, -76, -128, 117, -62, -124, -112, 12, 11, -9, 81, -78, 120, 102, -119, -56, 54, -69, 106, 10, -116, -1, 91, 32, 3, 22, 67, 101, 7, -68, -25, -24, -33, 61, 4, 64, 80, 81, -41, 63, -17, -101, -35, -59, -51, 120, -14, -61, -113, -15, -38, -10, 100, 64, 33, 46, -16, 26, -31, 22, 51, 52, -28, 53, 5, -66, 2, -41, -22, -13, 29, 109, 35, 6, -90, 71, -81, 26, -84, -111, 5, 2, 85, 125, 51, -81, -24, -39, 11, 11, -87, 101, 56, -59, 61, -119, -18, -74, 102, -124, -14, -3, -117, 8, -39, -121, 38, 36, 10, 111, -63, -101, -127, 45, -69, -105, -2, -84, 87, -126, 2, -59, 124, 66, -78, -112, 101, -48, -81, -53, -82, -52, 33, -35, -70, -95, -68, 8, -123, -87, 76, 33, -3, -105, 107, 13, 77, 117, -123, -127, -19, 11, -79, 55, -120, -120, 24, -73, 104, -25, 114, 65, -18, -18, -88, -122, 56, 91, 17, -128, 58, 43, -3, -60, 22, 20, 30, 46, 88, -73, -10, 38, 105, 45, 23, 45, -33, -37, -5, -46, -16, -1, -31, 76, 58, -52, -125, -23, 35, -35, 3, 116, 119, -43, -116, 105, -108, 53, 68, 114, -31, 91, -109, -95, 104, 89, -84, 23, -4, 57, -30, -96, 67, -48, -119, 28, 118, -120, -100, -117, 60, -73, -11, 102, -2, 120, 111, -37, -36, -110, -81, -83, 106, -75, -6, -55, 80, 35, 92, 32, 69, 16, -20, 88, 74, -43, -87, -62, 58, 118, 52, -104, 102, -121, 5, 86, 2, 104, 28, -104, 94, -63, 121, -87, 110, -118, 79, -18, 119, -15, 65, -62, -124, 4, -66, 55, -94, -51, 74, 77, 35, 14, 31, 103, 65, -19, -15, -64, -14, -62, -48, 17, -67, 58, -113, 78, 22, 94, 46, 73, -8, 23, -91, -104, 37, 69, 34, 87, -1, 115, 47, -14, -90, 121, 96, 11, -91, 84, 93, 87, -80, -112, 71, -123, -103, 13, -25, -127, 35, -122, -98, 120, 38, 86, -126, 109, 69, 79, 39, 50, -15, -126, 77, 113, -104, -117, 27, 31, -119, -88, -72, 10, 76, 0, 76, 105, -110, -56, -41, -119, -83, 106, -50, 49, -18, -48, -13, 55, 15, -39, 119, 118, -76, -29, -61, 109, -8, -31, 20, 77, -39, -67, 56, -110, -27, -28, -126, 44, -107, 39, 27, -23, -83, 23, 4, 46, 71, 90, -10, 89, 64, 77, -76, 18, -51, -15, 37, -67, -74, -39, -74, 49, 9, 92, -15, 3, -10, -94, -15, -44, 32, -50, 86, -18, -85, 55, -88, 32, -99, -79, -11, -31, 98, -11, 105, -73, 83, 10, -37, 20, -50, -51, 60, -29, 88, 81, -61, 90, -86, -2, -40, 13, 60, 116, 73, 111, 0, 25, -6, 95, 47, 111, 35, 12, -117, 98, -2, 100, 38, 123, -32, -26, 109, 64, -49, 125, -119, 94, -38, -68, 98, 91, 17, -37, 40, 107, -58, -69, -60, -36, 40, 123, -107, -92, -68, 18, -19, -35, -48, -5, 122, 10, -122, -25, 91, -114, 49, -124, 31, 27, -70, 65, -81, 112, 58, -45, 9, -30, 35, -27, -38, -20, 81, 15, 54, -12, 51, -47, -93, -20, -10, -91, 24, -27, -78, -5, -91, -81, -22, 57, 42, -40, -122, -48, 71, 75, 2, -114, 41, 109, 61, 113, 89, -97, -41, 59, 48, -107, -128, -127, 65, -5, 75, 108, 71, -85, -3, -39, -17, -29, -113, -120, 49, 38, -23, -106, 94, -118, 118, -32, 67, -104, 117, 76, -118, -26, 94, -67, -65, 65, 111, 88, 38, 112, 104, 73, 31, -9, -47, -48, 57, -37, -21, 71, -26, -60, 30, 64, 61, 109, -71, 127, 17, 35, 123, 126, -71, -91, 24, -14, 73, 28, -91, 127, 127, 26, -105, 113, -37, -90, -103, -90, 67, 0, 114, -118, 3, 87, -93, -33, 46, -39, 14, -114, -38, 31, 11, 124, -94, 59, 113, 9, 123, -57, -52, 91, -58, -84, 71, -8, 105, -46, -116, -119, 76, 38, -45, 107, -72, -120, 56, 21, -91, -38, 29, -99, 42, 16, 24, 114, 125, 22, 120, 25, -121, 39, 125, 99, -60, -2, -125, 112, -24, 23, -24, 112, 17, -104, 65, -116, 7, 5, 99, -12, -57, 102, 64, -117, -26, -48, 44, 4, 14, 32, -68, 92, 82, 81, -95, -67, 91, -116, -116, -92, -8, 40, -55, -72, -15, 80, -63, -86, 114, -115, 18, -89, -52, 108, -91, -65, 98, -29, 17, -104, 5, 85, -31, -85, 49, 52, -117, -94, 37, -45, 82, 0, -94, -106, 69, 0, -116, 7, -75, 2, 39, 74, -65, 78, -58, 69, 80, -90, -109, 49, 121, 18, -76, -65, 24, -65, 73, 13, 97, -63, -70, -82, 74, -115, -112, -65, -48, 2, -116, 121, 43, 39, 107, 91, -47, -5, 6, 66, 53, -6, 12, 98, 4, 88, -105, 103, 83, 110, -112, -88, 37, 11, -64, -98, 41, 120, -7, -49, -100, -6, -106, 64, -38, -92, -45, 62, 89, -28, -42, 14, 8, 93, 121, -1, -100, 64, -125, 39, -58, -117, 26, 36, -41, -118, -55, 100, -54, 125, -99, -22, -46, 110, 79, 26, 86, -115, 113, -61, 87, 85, 95, -30, 77, 60, -33, -16, 83, 8, 20, -114, 22, 82, 53, 57, 90, -128, 1, 55, -99, -77, 50, -54, 2, 121, -115, -122, 52, -6, 55, -96, 97, -33, -68, 63, 0, -8, -77, -23, 110, -63, 99, 23, -19, 35, -66, -105, -122, -22, -51, -115, 41, -98, 96, -16, -22, 13, 8, 97, -44, -122, 5, -5, -44, -19, -29, -83, -22, 67, -70, 59, -125, 90, 88, -53, 37, -66, -113, 94, 29, 16, -19, -115, -14, 73, -123, 123, -48, -6, -114, -21, 79, -81, 9, -112, 100, -3, -25, 57, -28, -3, 7, -11, -57, 62, -110, -44, 57, 69, -78, 48, 77, 119, -121, -3, -71, 100, 0, -108, 61, 38, 15, 90, -51, 52, -112, -62, 83, 127, 100, -84, -66, -19, 3, 119, 81, -8, 53, 34, 59, 100, 77, -22, 114, 78, -83, -23, -61, 67, -6, -101, 13, -94, 90, 76, 78, -39, 100, 32, -49, 81, -22, 15, -81, -104, 9, 53, 41, -8, -92, -124, -38, -91, -121, 43, 5, 82, -26, -15, 21, 70, 5, 126, 59, -104, 126, 63, 106, -100, 20, -77, -71, 20, -10, 100, -46, 73, -67, 80, 78, -54, 106, -12, -67, -75, 5, -70, -62, -91, -84, -22, 74, -39, 127, -117, 9, 17, -45, -7, -105, -15, 23, 32, -44, 124, 8, 94, -41, 72, -79, 96, 20, 47, 123, -50, 86, 16, -128, 49, 98, -92, 91, -39, -21, 84, -73, -85, -47, 39, 18, -14, -115, -27, 7, 92, 54, -53, -127, -54, 80, 28, -27, -54, 32, -54, -28, -100, -83, 106, 29, -30, 32, 89, -107, -52, -103, 80, -125, 124, -78, 16, 89, 26, -1, 15, 47, -121, -31, -70, -14, -22, -114, 51, 67, 117, 83, -9, -6, -110, 60, -64, 25, -60, 95, 89, 65, 89, 11, -112, -105, 127, -123, 114, -24, 52, 56, 103, -3, 7, 70, -68, 32, 107, 43, 45, 41, -27, 78, -52, 121, -17, 125, -34, -52, 37, -7, 46, -92, 47, 77, 59, 94, -76, -63, 27, 4, 109, 101, -19, -24, 39, -27, 93, -122, -119, 31, -58, -111, -44, -76, -30, 23, 25, -126, 34, -80, -35, 56, -101, 4, 120, -113, 97, 74, 43, -98, -26, -112, -65, 108, 41, 113, 124, -45, 11, -5, -77, 70, -13, -15, -14, -20, -46, 85, 120, 88, 0, 20, 70, -51, 111, -90, -25, 116, -1, 111, 100, -106, -71, 78, 117, 31, 89, -1, 0, -69, 34, 88, 3, 22, -127, -92, 112, -124, 73, -27, -7, -80, -105, 54, 82, 116, -48, 75, 76, 40, -13, 113, 35, 47, -124, -114, 107, 38, -47, 86, -95, -101, 90, -15, 90, 48, -42, 59, -120, -95, -32, 69, -105, 120, 102, 96, -63, -124, 87, 119, 8, -72, -99, 9, -90, -55, -97, 114, 107, 100, 99, -79, 59, -86, 40, 90, -81, 31, -82, -114, -78, 10, -80, 108, -87, -55, 93, 115, 80, -38, 70, -99, -110, -98, 65, -89, 105, 25, 67, -33, 29, -9, -99, 113, -57, -23, -24, -96, -121, 74, 97, -32, 11, 1, 24, 112, 123, 43, -30, 117, 15, -50, -22, -85, -13, -111, -128, 95, -49, 11, 78, -120, -16, 53, -106, 17, 91, 12, 6, 112, -95, 11, 107, -17, -32, 12, 58, 123, -124, -72, 67, -37, -85, -17, 67, -82, -109, -125, -113, 16, -75, 107, 29, 124, 84, 67, 98, -69, -12, 99, 45, 105, 120, -96, 69, 11, 42, -33, 18, 62, 65, 71, 107, 15, -67, 99, 12, 69, -66, -103, -91, 30, 75, 61, -115, -75, -63, 16, -93, -91, 1, 77, -20, 61, 20, 108, 109, -79, 62, 54, -29, -61, 80, -72, 79, 75, 36, 39, 8, 53, -83, 60, 37, -6, 3, 73, 20, -2, 28, 52, 63, -100, -120, -32, 82, -48, -14, 49, -64, 53, 73, -50, 116, -36, -123, -106, 37, 23, -27, -113, -83, 98, 86, 20, 94, -115, -82, 7, 35, 30, 64, 40, 112, 48, 95, -18, 103, -126, 7, -36, -101, 72, 107, 56, -52, 60, 106, 64, 73, -28, -106, -1, 57, 73, 104, 33, -34, 2, -42, 31, 6, 110, 33, 127, 123, 88, -32, 50, 15, 76, 61, -126, -110, 26, 39, 54, 17, -27, -55, -56, -57, 122, -35, -9, 70, -37, -72, -26, -102, -77, 7, -121, -76, 119, -111, 38, 88, 39, -1, 15, -96, -37, 127, -81, -14, -109, 120, 119, -21, -46, 121, 45, -60, -10, -28, 56, -24, 122, 15, 109, -43, -71, -91, -57, 94, -15, -127, 127, 65, 11, -119, 54, 97, -40, -72, -36, -9, -85, -80, 7, -128, 81, -119, -36, -41, -115, 77, -55, 103, -43, 6, -88, -84, 64, 1, 95, -118, 112, 106, -77, -3, -30, -22, 110, -71, -15, 65, -71, -33, -32, 127, -22, -127, 61, -53, 112, -80, 78, -91, 101, -76, 17, 60, -77, -25, -64, 50, -18, 85, 109, 79, 75, -44, -78, 97, 77, -66, 36, -7, 15, -56, -91, 92, -125, 6, 41, 45, -12, 86, 40, 25, 43, -43, -100, 68, 56, -106, -61, -73, 26, 83, 90, -5, -118, -20, -10, -13, 12, 53, 106, 105, -98, 67, 37, 32, -40, -111, 23, -42, 107, 34, -110, -69, 74, -108, 88, -5, 41, -55, -80, -62, -112, -19, 27, -100, 1, 103, 64, -84, -68, 51, 65, 118, 114, 104, 7, 80, 74, 26, 96, 19, -58, 64, -7, -85, 103, 54, 17, -79, 49, -113, -56, 112, 127, 104, -106, -122, 58, -11, -120, -41, -117, -32, -6, -104, 86, 68, -57, 46, 114, 93, 74, -119, -69, -20, 13, 103, -18, -21, 42, -85, -4, 36, -44, -93, -103, -47, -17, -18, -119, -47, 89, 117, -23, -35, -122, -114, 31, -10, 10, -34, 30, 23, -116, -105, 27, 106, 40, -109, 42, 38, -83, 98, 79, -128, -9, -27, 13, -11, 7, -50, -86, -50, 93, -27, 56, 89, -29, -16, -84, -53, 111, -109, 95, -104, 21, 62, 107, 31, 45, -82, 33, -11, -27, -25, -41, -87, 119, -110, -33, 55, 69, 22, -62, -28, 95, -91, 105, -63, -122, 111, 19, 65, -49, -73, -75, -8, 71, -22, -57, -15, -94, 44, -22, -61, 31, 7, -39, 126, -108, -63, -29, 114, -56, -91, -70, -11, -9, 42, -95, -25, -42, -116, -95, -55, 69, 77, -54, -32, -110, -33, -26, 126, 125, 108, -89, -42, 70, 36, -111, -127, 40, -84, 118, 24, 64, -21, 79, -95, 86, -14, -78, 70, -59, 61, -88, -87, -37, 113, -69, -102, -37, -56, -89, 38, 75, -27, 12, 104, -109, -55, -111, -51, -96, -102, -57, -47, 48, 32, 9, -104, 42, 59, -2, 58, 24, 39, -16, 102, -26, -72, -42, 117, -128, 62, -23, 9, -124, 30, 66, -126, -58, -70, -93, -128, -7, 60, 73, 116, -35, 56, -84, -108, -89, -22, 77, 77, -125, -100, -17, 105, -112, 58, -57, 73, -101, 74, -2, -80, -55, -41, -26, -69, 74, 80, -75, 47, 3, -94, -50, 126, -70, -30, -28, -111, -15, -42, 81, -2, 108, 44, 51, 65, 35, 121, -107, -84, 47, -72, -17, 79, 29, -42, -60, 120, 104, -34, -98, 42, 31, -62, -26, 39, -96, -127, -37, 89, 32, -58, 116, -69, -27, -11, 68, 34, 53, 25, -93, 88, 34, -54, 52, 44, -104, -70, -14, 19, 72, 118, -120, -46, 29, -125, 83, 14, 79, -3, 87, -81, -110, 104, 25, 97, -107, -31, 52, -88, 45, -122, 78, 12, 27, 99, -78, 124, -70, 121, 19, 111, 18, -31, 15, 70, 56, 126, -98, 69, 23, -83, -52, 127, -15, 50, -60, 55, 39, -113, 19, 115, -32, 98, -64, -2, 25, 14, -9, 0, -103, 60, -37, 75, -25, -52, 22, -72, -15, 12, 94, -86, -7, 107, 4, 64, 20, 86, 124, -103, 93, 66, 110, -95, -49, -116, 8, -107, 110, -10, 32, 66, 83, -48, -121, -44, 65, -66, -121, -65, -15, -99, -71, 54, -92, -25, -117, 56, -42, 94, 107, -69, -101, -57, 122, -41, 95, -18, -15, 95, -42, 10, 18, -3, -78, 84, 81, -13, -30, -18, 77, 69, 20, 21, 20, 49, 83, -5, -90, 48, -62, -85, 26, -57, 124, 86, 22, 0, 3, -23, -59, -3, -95, 48, 108, -25, -85, 18, 28, 117, 37, 125, -70, 108, -76, -100, 13, 93, 107, 43, 6, -40, 3, 98, -57, -51, 53, -128, 4, 125, -3, 57, 105, -110, 112, 123, 58, -15, -18, 73, -101, 58, 16, -54, -35, 87, -110, -80, -84, -10, 1, -116, 16, 28, -41, -120, 110, 27, -37, 58, -21, -51, -104, 64, -97, 28, -65, 77, -98, 112, -96, 108, 27, 40, 80, -53, 116, 50, -67, 25, -85, 16, 20, 60, -47, 12, -32, 88, -57, -22, -83, -59, 53, 98, 91, 67, 45, 51, -8, 19, 20, 12, 114, -12, 66, -59, -28, -38, 39, 95, 2, 126, 102, -62, -96, -101, 59, 7, -91, -53, -8, 40, 111, 96, 90, -128, -123, -25, 97, 118, 80, 86, 20, 30, -112, 14, -125, -30, -32, 122, -114, 35, 115, -73, -32, 36, 65, 101, -27, -79, 7, -122, 9, 83, -119, 54, 32, 90, 77, 11, 75, 4, 10, 25, 111, 73, -8, 127, -41, 11, 113, -24, 6, -38, -38, -106, -88, -12, 114, 114, -102, 112, -92, 65, 11, -12, 17, 86, -6, -33, 3, -57, -93, 21, 38, -4, 10, -28, -39, -16, -62, 126, 88, 29, 28, -106, -25, -47, 101, -7, 20, -60, -56, -63, 50, -73, -127, -60, 28, -113, 30, 114, -94, -2, -49, -39, 1, -28, 15, -118, 43, -98, 14, 5, -9, -113, -100, -42, 86, -80, 51, -28, 50, -47, 40, 50, -1, 77, -120, -109, 72, -91, -112, -100, 26, 30, -86, 122, -20, -96, 63, 41, 48, -100, -8, -2, 98, 90, -101, 83, 50, 84, 104, -81, -74, 24, -78, 34, 95, -12, 50, 5, -106, 47, 96, 81, 112, -117, 108, -112, -50, 28, 126, -47, -38, -90, 57, -7, -82, -112, 82, 67, 114, 118, -83, -27, -6, 122, -115, 119, -9, -2, -52, -27, 65, 9, -113, -23, -86, 10, 88, -59, 58, 47, -23, 112, -81, -57, -24, -15, -120, -83, -79, -91, -4, 96, -41, 2, 65, -95, -101, -49, -76, 111, 78, 21, -33, -62, -95, -7, 104, -54, -102, 69, -46, 17, 115, 14, -88, -37, 22, -87, 63, 48, -17, -108, 21, -109, 100, -68, -34, 116, 66, 3, 59, -97, 94, 50, 82, 127, 92, 80, -95, -54, -107, 113, 87, -26, -55, 103, -68, -3, -18, 32, 46, 63, -24, -113, -63, -81, -56, -98, 127, 65, 122, 13, -81, -121, -77, 108, -39, 45, 12, 53, -65, -14, -116, -96, 8, 14, 7, -110, 52, 125, 28, -69, 103, 35, 105, 0, 29, 109, -69, -82, 29, 30, 102, -71, 36, -76, 81, -77, -35, 7, 122, 56, -93, 60, 116, -10, -127, 17, -53, -64, -62, -108, 23, -91, -92, 91, -107, -111, 40, -72, 40, 2, -99, -78, -70, -7, -6, 18, -73, 78, 69, 57, -84, -55, -116, 59, 14, -102, 117, -110, 40, 118, -123, -50, -33, 123, 97, -93, -87, -80, -32, 110, -78, 92, -95, 123, -95, -39, -61, -12, 33, 41, 36, 9, -40, 28, 13, 28, -18, -55, 43, -50, 3, -33, -23, -20, 56, -91, -100, 0, 25, 48, -107, 113, -78, 102, 79, -6, 68, 72, 102, -33, 12, 79, -104, -6, -21, 17, 101, 123, -114, 53, 127, -128, 120, 111, -125, 1, 114, 64, 42, 119, 81, 48, -49, -128, -105, 7, -40, 96, 87, 98, -28, -18, 84, -96, -109, -94, -61, -61, 124, -99, -106, 84, 60, -59, -13, 30, -46, 81, 35, 38, -71, 71, 91, 82, -44, 74, -4, 92, 124, -9, -116, -39, 18, 24, 6, 29, -32, -117, 15, -76, 43, 23, 11, -120, 73, 1, -69, -54, 64, 18, -22, 100, 85, 49, -54, -75, -51, 120, -108, -78, 71, 90, -27, 97, -110, -24, -69, 51, -83, -102, -56, -48, -19, 91, -52, -95, -18, -112, 60, 59, -33, 126, 73, 44, -96, 114, 3, -122, 83, 32, -62, -126, -3, -27, 119, -58, -114, -99, -65, -93, 54, 109, -24, 28, 55, 60, 40, 46, -91, -56, 112, -118, 87, -50, 104, -29, -34, 123, 123, 97, 47, -108, -114, -50, -94, 70, -96, 3, -73, 126, -54, 94, 78, 40, -82, 30, 70, 91, 118, 68, -10, -78, -12, -1, -8, 75, 98, -22, -62, -123, 98, 84, 66, 122, -106, 60, 81, 92, -47, 13, -94, -34, 59, 118, -107, -63, 89, 43, 65, -55, 63, -123, -90, 108, -85, 59, -24, -19, 13, -8, -74, 104, -118, -118, 12, -74, -67, -44, -24, 94, 93, -111, -113, -98, -21, -80, 10, -89, -60, -108, -13, -27, 48, 14, 22, -31, 95, -107, -126, 107, 32, 11, 5, 20, -82, 108, 44, 94, -79, 106, -9, 73, 80, 87, 47, -27, -34, 77, -93, -94, 95, 87, -112, 39, -72, -56, 74, 19, 6, 35, -105, -15, 106, -90, -91, -3, 13, 116, -97, 69, 3, 101, 65, -39, 73, -29, -22, -24, 90, -62, 16, 116, 40, -115, -25, -4, 15, -19, -37, -32, -42, -24, 42, 45, -125, 51, -119, -74, 80, -68, 115, 91, -20, -71, 19, 75, 86, 77, -67, -12, 8, 14, -28, 87, 25, -40, 87, -14, -57, -5, -115, 27, 91, -93, -67, -67, -120, -47, -65, -78, 24, -72, 74, 74, 90, -118, 106, 103, 111, 74, 115, -27, -128, 46, 34, 80, 77, -122, 33, 124, -77, 9, -63, -75, 59, 112, 20, -37, -47, -35, -94, 63, 110, -95, 110, 27, 52, 47, 71, 3, 45, 33, 115, -46, -90, -35, 53, -7, -11, -62, 91, 43, -14, -68, -121, 30, 23, -1, 58, 106, 84, -9, -119, 59, -91, 6, -49, 2, -51, 63, 61, -22, 89, -104, 127, -92, -26, 15, -79, 24, 111, -11, 108, -112, 3, 66, -97, -103, 64, 116, 17, -35, 42, 71, 11, -84, -100, 78, 15, 89, 105, 74, 94, -40, -4, 119, -82, 37, -2, -52, -31, 45, -67, 59, -1, -117, 8, 77, 55, -91, -71, 29, -62, 2, 103, -107, -2, 99, -42, 74, 39, -96, -44, -44, -108, 92, -55, -53, -110, -120, 92, -56, 17, -44, -112, 16, 41, 75, 96, -104, -101, 97, -10, -72, 116, 15, -101, -85, 70, 43, 56, 80, 76, -29, -92, 124, 119, 8, -108, -40, -91, -84, 81, 119, 21, -43, 0, 82, -102, -60, -122, 49, -30, -70, 78, 17, -13, 100, 58, -60, 6, 92, 2, 28, -21, -115, -9, 77, -50, 75, -56, -110, 5, -126, -39, 0, 60, -115, 10, 14, 64, 93, -75, 94, -104, -71, 3, -101, -55, 15, 122, 31, 19, -63, -128, 115, -95, -9, 0, -90, 94, -15, 115, -64, -36, 23, 87, -52, -102, -111, 81, -39, -76, 3, 76, 95, -34, -3, -108, 103, -4, 37, -13, 88, 4, 37, 114, -97, -83, 66, -100, -55, -123, 37, -82, -105, -31, -102, 92, 84, 110, -35, -80, -58, -48, -2, 35, -80, 100, 80, 102, 84, -48, 7, 10, 37, -15, 5, 97, 13, 8, 75, -122, -84, 102, 51, -121, -73, 10, 84, 12, -122, 119, -116, -61, 123, 69, 95, 123, 1, 16, -24, 20, 59, 30, 102, -77, -58, -27, -63, 103, -58, 127, 10, 27, 69, -107, 44, -126, 51, -56, -74, 104, -127, 79, 63, -102, -8, 114, -62, 107, 127, 91, 18, -21, -43, -112, 125, -71, -25, -109, -6, -118, -36, -64, 4, -109, -26, -13, 28, -91, -63, -56, 41, 7, 52, 0, 35, -9, -63, 74, -56, -68, -38, -66, 43, 55, 105, 83, 105, -44, -50, -42, 41, -107, -124, 98, -114, -31, -111, -104, -9, -36, 98, -121, -16, -110, 67, 47, 74, -78, -82, 64, -121, -113, -118, -94, 69, -91, 70, 15, 27, 58, 11, -96, -115, 66, 85, -47, 48, -34, -121, -52, 31, -104, 6, 118, -3, 51, 54, -34, 108, -9, -49, -60, -7, -125, 40, -80, 40, -123, 41, 45, -101, -14, 43, 100, -68, 5, -123, 70, 125, -81, -62, 40, -47, 0, 122, 103, -27, 52, -120, 94, -95, -70, 74, 58, 0, -39, 61, 40, 88, -103, 79, 5, 6, 103, 26, -55, 27, -81, 43, 71, -86, 47, 120, 48, -121, 41, -16, -62, 12, -43, 66, 74, -98, 113, 121, 122, 63, -105, 50, -95, -6, -59, -73, 44, -75, -89, 74, -70, -80, 26, 59, 53, -37, 80, 9, -47, 108, 123, 46, 30, 49, 72, -35, -5, -67, 82, 115, 102, -46, -51, 3, -58, -61, 71, 49, 62, 93, -25, 59, 56, -29, -70, 31, 21, 83, -127, -76, -56, 28, 30, -115, 72, -30, -4, -104, 13, 67, -15, 125, 77, -24, 11, -42, -56, 95, 53, -84, -31, -15, -81, -110, 52, -72, -22, 102, -127, -80, 95, -93, -9, -120, 81, -4, -56, -123, -87, 5, 50, 108, -64, 54, 116, 98, 120, 13, -52, -5, 119, 43, -118, -17, -23, -34, 7, 100, -91, -100, -30, 64, 83, 92, -75, -55, -53, 118, -30, -75, -128, -9, -20, 66, 59, 88, 90, 119, 5, 113, 50, 5, 109, -114, -124, 27, -45, 120, 4, -41, -100, -37, -100, 37, -111, -28, 115, -111, -79, -1, -124, 84, 46, -85, 73, 1, 89, 20, -99, 18, -15, 125, 82, 56, -1, -62, -18, 59, 69, -24, -75, -87, -81, 27, -87, -59, -51, 74, -44, -118, 47, 30, 124, -105, 81, -5, -71, -72, -17, 100, -70, -39, -54, -34, -85, -14, 68, 107, -77, -38, 37, 38, 121, -73, 121, -77, -2, 52, 108, 117, -8, 31, -75, 71, -106, 47, -42, 107, -67, -126, 4, -10, -34, 55, 21, 4, -85, -120, 43, 11, -92, 43, 63, 59, -18, -56, -37, -73, -115, -1, -26, -9, 60, 31, -29, 126, 55, -70, 117, -65, 112, -86, 122, -101, -92, 64, 16, -111, 108, -32, -71, -39, -110, 44, 21, 57, -77, -47, -69, -83, -6, -49, -14, 76, -10, -56, 86, 90, -50, -20, -103, -64, 113, -28, 24, 65, 80, -39, 114, 38, 93, 31, -31, 118, -70, -64, 15, -103, -81, 87, 60, -28, -76, -90, 98, 10, -50, -2, -36, -80, 41, -26, 33, 41, 33, -122, -10, -52, 41, -91, -3, -118, -117, -91, -105, -12, 125, 87, 117, -103, 24, 119, -57, 110, -65, 124, 9, 51, -42, 78, 30, -113, -89, -123, 30, -23, -76, -36, -82, -7, 71, 36, -96, -113, -16, -95, -27, 101, 95, 88, -123, -57, 112, 37, -122, -52, 43, 120, 12, 75, 32, 110, -118, 103, 65, 34, 102, -104, -103, 8, 88, 93, 105, -97, 98, -21, -73, 120, 86, -127, 41, -58, -110, -97, 119, -92, -100, 122, 117, 16, -5, 31, -117, 47, -117, 83, 127, 15, 88, 94, -60, 2, -25, -14, -118, -116, -116, -47, 26, -6, 63, -117, -127, -68, 92, -50, -59, -23, 101, 109, -45, -32, -12, 2, 57, -84, -6, 2, -57, 76, -24, -121, -40, 18, -23, -4, -119, -53, 107, -65, 61, 91, -59, -22, 97, -36, 0, -101, -91, 68, -126, -78, -93, 55, -96, 96, -7, -86, -99, 54, 39, -96, 126, 67, 79, 15, 75, 103, 49, -48, -12, 102, 67, -104, 82, -11, 39, -107, -74, -79, 31, -19, -104, -110, -2, 0, -82, 12, -74, -63, -114, 117, -51, -102, 63, 114, 0, -39, -56, 23, -96, -63, 34, -47, -76, 76, -71, 76, 121, -90, -74, 92, 67, 18, 22, -97, 25, 38, 39, 77, 51, 76, -42, -120, -10, 94, 89, 95, -69, 57, -59, -112, 42, 60, 57, -42, -68, 119, 28, -36, 118, -124, -114, 120, -97, -81, -23, -23, 79, 110, 23, -14, -122, -25, -73, -99, 88, 70, -4, -69, -91, 118, 120, 28, -62, 49, -16, -94, -123, 126, 47, 124, 67, -70, 86, 22, -55, -42, 89, -115, -16, 104, 35, 113, 124, 88, -54, 75, 5, 61, 3, -1, 19, -86, -70, 34, 100, -49, -125, -19, 9, 100, 111, -78, -12, -41, -81, 120, 124, 127, 122, -76, -84, -47, 52, 16, 124, 2, -125, 40, 7, -22, -11, -120, 22, -68, 49, 109, 101, 116, -107, -126, -96, 96, -125, -73, -64, -3, -38, -6, -36, 20, 21, 51, 107, -102, -20, -23, 0, 31, 0, 10, -90, 103, -71, -21, 67, -59, -41, 79, 43, -51, -100, -124, 14, 14, 24, 43, 77, 123, 38, -17, -92, 38, 80, 27, 50, 18, -83, -99, -108, 97, 99, 80, 91, 85, -61, -80, 45, -114, 0, -104, 127, -40, -69, 126, -93, -2, 111, -65, 54, -82, 14, -19, -92, -96, -93, 34, -105, -57, 9, -26, 18, -28, 32, 87, -44, -76, -24, 61, -43, -88, -21, 79, -38, -5, 103, -97, 78, 99, 77, -115, 110, 100, -30, 18, 23, -101, -77, -95, -72, 119, -53, -55, -21, 90, -101, -76, -121, 23, -29, -90, -47, -10, 24, 15, 4, -40, -1, -70, -121, -65, -4, -47, 24, 11, -17, 15, -99, -45, 24, -90, 33, -36, 7, 52, 76, -104, 89, 90, -12, 6, 72, -108, -21, 97, -119, 118, -28, -123, 101, -37, 22, 127, -67, -30, 75, -47, 43, -125, 95, 25, -116, 27, -127, -53, -32, 86, 14, -121, 111, 10, -126, 71, -4, 109, 81, 98, 4, -38, -4, 70, -110, 98, 47, -99, 88, -114, -127, 99, -83, -53, 66, -34, -75, 67, 54, -71, 84, -13, -81, -8, 82, 60, -126, -38, -74, -76, 12, 31, -9, -92, 122, 122, -31, -66, -99, 114, 63, 86, 80, 72, -38, 84, -102, -40, -87, -39, -9, -108, 29, 71, -86, -20, -113, -120, 72, -57, 80, 94, -47, 89, 6, -21, 35, 65, -115, 53, 38, 40, -24, -98, 26, -37, 33, -7, 97, -7, 114, -37, -83, -47, 63, 35, 14, -112, -99, -51, 57, 122, 93, -57, -88, -4, 114, -35, 3, 79, -49, 100, -120, 88, -42, 98, 37, 106, 106, 33, -19, -111, -74, 108, 47, -57, -83, 89, 78, -2, 83, 66, 86, -66, 116, -114, -36, -60, 43, 46, 3, 5, -104, 20, -102, -50, -70, 40, -45, 32, 92, 93, -105, 120, -87, 59, -20, 85, -96, -51, 122, -81, 53, -17, -120, 16, -27, -64, 11, 35, 52, 116, 119, 122, 12, 51, 109, -26, -70, 78, 98, 99, -33, -29, -71, -14, 90, -78, -82, 77, 38, 100, 123, -109, -45, -1, -11, -82, -33, 111, 38, 21, -29, -40, 73, -45, 66, -92, 111, -48, -89, 31, -117, 79, -27, 36, -85, -49, 6, 55, 97, 54, 4, -36, 23, 68, -18, -47, -105, -34, -62, 81, 2, -14, -69, 33, 69, -43, 124, 17, 99, 107, -6, 60, 98, -92, 15, 112, 115, -73, -72, 110, 58, 99, 115, 4, 50, -39, 106, -32, 75, -55, 50, -17, -108, 102, -31, -18, 79, -43, -87, 17, 10, 16, -111, 21, -82, 19, 44, -67, 2, -111, -23, 25, 7, -19, 65, -110, 52, -60, -63, 102, 106, 27, 89, -87, 104, -38, 43, -114, 2, -49, 78, 111, -11, -13, 18, 10, 3, 120, -43, 88, 114, -110, -50, -89, -44, 76, 65, -16, -123, -106, 68, 49, -41, 107, 64, -111, -66, -4, 55, 21, 86, 2, -107, 115, 99, -89, -58, -112, 116, -127, 44, -21, 83, -128, 54, 7, 41, 12, -90, 79, -67, -89, 61, 35, 90, -21, -58, 69, 5, -13, 51, 71, 61, 25, -106, -22, -105, 86, 60, -33, 48, -9, 108, 5, 56, 41, -38, -94, -70, 22, -76, 3, 19, 42, 41, 47, 37, 80, -74, 48, 30, 127, -123, 52, -85, -5, -7, -69, -105, -99, 99, 84, 66, 42, 46, -123, 58, 69, 62, -88, 62, 122, -124, 75, -102, -85, -45, 81, 123, 33, 82, -114, 25, -90, 69, 105, -20, 120, -76, 60, 40, 10, -123, 60, -116, 26, -70, -58, -102, -65, 6, 35, -55, -103, 33, -45, -102, 33, 28, -123, 5, -18, -87, -32, -9, 28, -18, -117, 38, -20, -48, 111, 7, -111, 56, 28, 62, -1, -42, 64, -79, 67, -58, 88, 68, -75, 22, 60, -108, 104, 41, 14, 73, 105, 32, 22, -52, 35, -79, -100, 90, 33, -94, -59, -75, -37, 74, 99, -33, -38, -100, 47, -92, 66, 103, 118, -67, -95, 12, 54, 11, 91, -106, -38, 37, -18, 57, -117, -27, -102, -67, -31, 117, 76, -92, -117, 31, -122, 116, -44, -93, 45, 66, 95, -59, 92, 82, 86, -78, -19, -94, -75, 11, -77, 105, 48, -125, 78, -69, -102, -96, 15, 16, 30, -79, 84, -62, 40, 118, -96, -5, -83, 121, -92, 14, 51, 34, 96, 123, 105, -72, 36, 82, 57, -55, -58, -25, -127, 123, 34, -128, -89, -39, -71, 120, -69, -29, 18, 87, -97, 41, -76, 50, -26, 97, -98, -109, 78, -98, -54, 105, -42, 48, -78, 56, -54, -81, 119, 10, -40, 0, 63, 15, 110, -93, -66, 122, 124, 65, -9, -45, 116, 76, 80, -1, 17, 3, 113, 120, 107, -88, -94, -76, 50, 97, -6, 29, 72, 1, -1, -93, 88, -124, 99, 8, 23, 52, -3, 18, -84, -36, 48, -17, -40, -109, -9, -78, -104, 30, -124, 35, 52, -59, 41, 95, -1, 72, 96, -109, -128, -8, 69, -38, -95, 81, 121, -70, -63, -38, 80, -98, -49, -57, -54, 118, -46, -54, -19, -115, -92, -120, 55, 42, 41, -16, -76, 17, 5, -31, -83, -87, -94, -110, 95, 75, -85, 17, -75, -7, 67, -27, -2, -8, -56, 111, -103, -111, -68, -38, -53, 19, -68, 73, -66, 25, 123, 18, 64, 22, -93, -5, -18, -93, -65, 54, -15, 116, -12, 65, 24, -85, -54, -29, -9, 93, -60, -107, -14, -20, -125, -23, -11, 121, 56, 121, 25, -2, -6, -22, 5, 100, -39, 76, -27, 113, 115, 111, -18, 123, -59, 110, -98, 62, 110, 51, -6, -110, -13, 71, -40, -70, -63, 11, 91, -12, -98, -58, 64, 80, 72, -4, 100, 34, 7, 47, -9, 104, -101, 46, -92, -46, 62, -58, 9, 124, -113, -126, -72, -123, 26, -67, -47, -14, -53, 44, 100, 31, -104, -60, -97, -119, -100, -52, 60, 11, -85, -69, 7, 103, -83, -51, -112, -36, 0, -2, 36, -20, -88, -28, 26, -78, 121, -63, -114, 33, 60, 34, -55, -82, -98, 68, -108, -103, -75, -51, -55, 90, -37, 64, 13, 78, -41, 37, -73, 12, 94, 15, 94, 37, 109, -5, -65, 3, 87, 8, -90, -68, 81, 120, 75, -34, 51, 5, 82, 72, -43, -118, 23, -18, 127, 23, 4, 122, 77, 54, -2, 59, 74, -26, 18, 50, -8, 106, 107, 72, -87, 113, -103, -122, 111, 111, 47, -26, 41, -105, 99, 77, -99, -84, -71, 10, -41, -2, -86, 32, 25, -15, 58, -40, -88, -39, -6, -127, -102, -111, 2, 39, 124, 58, -88, 4, 30, -80, -119, 116, -63, 90, 109, 57, -6, -92, -88, -116, 76, -115, 125, -10, 17, -78, 119, 110, -21, 80, 120, 47, -112, 58, -122, 43, 107, -123, -107, -59, 56, -91, -6, -3, 71, -105, -66, 69, -29, -20, 51, 24, -34, 105, 61, -83, -31, 38, 26, 67, -122, 95, -103, -113, 49, -11, 80, -59, -110, 63, -89, -70, -78, -51, 34, -49, -4, 100, 104, 99, 45, 76, -111, 25, -101, -26, -80, -43, 108, 113, 121, 79, -107, -76, -123, 48, -77, 45, 30, 3, -43, 91, -42, 126, 18, 123, 80, 16, 108, 87, 126, -119, -73, -111, -40, 53, -65, -84, -31, 66, 100, -73, -4, 23, 33, 36, 89, -123, -89, -55, -62, 50, -74, -113, 17, 91, -59, 55, 30, 2, 15, -7, 26, -27, -33, 122, 77, -73, -95, -45, 115, -84, 30, -92, -90, -91, -101, -124, -83, 107, -125, 38, -5, 108, -35, 92, 73, -90, -50, 43, -74, -112, -97, -32, -84, -21, -16, -103, -37, 36, 66, -28, 0, -110, 98, -13, 11, -72, -126, -78, 95, -81, -44, -96, 90, 69, 71, -103, 8, 77, -88, 77, 36, 50, 68, -54, -16, -121, -114, -74, -95, -25, 57, -36, -67, 62, -6, 76, -39, -16, -32, 45, 95, -16, 13, -102, -8, -71, -12, -50, 34, 25, -6, -10, -114, -36, 66, -42, -116, -46, 103, 56, -14, 114, 45, 98, 89, 18, -108, 55, -67, 40, 108, 83, 105, 33, 105, -109, 31, 120, -81, 107, -119, 40, 95, 44, 56, 68, -105, 22, -80, 18, -35, 116, 93, 63, 51, 124, 96, 82, 123, 62, 125, 108, -33, 51, 77, -36, 57, -119, 52, 70, 64, 43, -64, -44, -108, 65, 73, -13, -125, 105, 127, -88, -41, 103, 79, -43, 15, 109, 125, -89, -127, -121, -87, -38, -41, 32, 32, -94, 91, 74, 95, 41, -20, -35, -61, 74, 75, 27, 70, 45, -20, -96, 17, 69, 52, -108, 8, -37, 119, -53, 41, -111, 108, -52, 16, -54, -34, 49, 17, -100, -107, 72, -110, -73, 84, -89, -47, -108, 20, -12, -42, 126, 37, -19, 60, -79, 36, 34, -70, -100, -64, 99, -83, 31, 2, 119, -21, 118, -127, 77, -102, 3, -17, -61, 95, 80, -96, -87, 61, 59, 90, -88, -105, 77, 12, 16, 24, -71, -114, -10, 22, -28, 124, 99, 120, -68, -91, -111, 114, 67, -27, 94, 2, -24, -84, -120, -23, -107, -38, 3, -52, 65, -14, -67, 28, -103, -126, -72, -15, -111, -68, 86, -106, -92, 40, 70, -40, -31, 96, -58, 0, 58, -66, -71, -28, -124, -5, -92, 19, 89, -102, 101, -119, 94, -88, 87, -62, 108, 106, -64, -108, -127, 76, -119, 80, 101, 119, 52, 76, -93, -128, -108, -13, 35, -20, -48, 41, -91, 81, -4, 116, -90, 121, -100, -100, -77, 23, 90, 56, -41, 111, 103, -48, 125, -24, 51, 110, 107, 96, 47, 79, 24, 67, -9, 68, -91, 82, 67, -100, 92, -17, 52, -16, -5, -2, 40, 26, -46, 108, 72, -86, -88, 82, -52, -84, 21, 4, 77, 59, -70, 27, -60, 84, -10, 43, -10, -51, 29, -14, -37, -99, 70, -32, 1, 52, -46, 122, 112, 51, 19, -67, -100, -78, 24, 118, -81, 5, 93, -114, 46, -47, -76, -86, 127, -34, 107, -49, -57, -114, 96, 119, 75, 45, 93, -61, 53, 2, 78, -9, -59, -38, 11, -52, 126, -118, -39, -111, 39, -52, 75, -25, -45, -116, -20, 93, -128, 23, -48, 0, 127, -118, 10, -34, 113, 25, -84, -40, -114, 88, 33, 34, -28, 102, 120, 73, 109, 18, -123, -53, -30, 11, 72, -68, -123, -66, -17, -26, 113, 38, -107, -101, 114, -12, -106, 127, 19, -22, -128, -27, -29, 92, 62, -76, 45, 97, 69, 48, 12, -8, -80, 71, 67, -78, -118, -91, -102, 88, 15, 100, -128, -23, -126, -77, 71, 62, 107, 11, -67, -84, -106, -75, 58, -25, -35, 55, 33, -65, -128, -42, 22, -102, -14, 26, 71, -30, 108, -1, 72, -36, -93, -45, -124, 43, 122, -105, -81, 4, 1, 102, -55, 68, -113, -24, -33, 34, -82, 123, -10, 48, 103, 78, 70, 50, 77, 34, 86, 62, 33, 37, 81, 76, 53, 20, -83, 75, 45, -60, 68, 72, 65, 93, 89, -6, -112, 43, 82, 94, 2, -22, -104, 12, 55, 50, 13, -39, -95, -70, 71, 23, 31, 39, -35, -9, 83, 9, 99, 14, 1, -38, -84, -115, -58, -3, 90, 6, -68, -124, 123, 90, 43, -80, -84, -84, 103, 32, 44, 70, 58, 56, 75, 117, -116, 106, 111, -119, 101, 89, 27, 109, -92, -17, -53, 47, -37, -43, 3, -50, 59, -43, 115, -128, 110, -80, -40, 113, 38, 107, -82, 17, 12, 2, 47, -8, -12, -24, -54, 112, -16, 78, -90, -109, -82, 60, 115, -43, 127, 33, -109, -88, -28, 102, 92, 91, 16, -53, -31, 89, -63, -45, 22, 27, -25, -69, -113, -116, 25, -112, 37, 69, 110, -66, 93, 60, 25, -66, 6, 57, -48, -10, -87, -51, 10, -65, 124, 100, 25, 58, -45, 64, 127, -113, -126, 59, 44, -95, -122, 91, 99, 92, -78, 3, -96, -93, -102, -73, 23, -42, 60, 89, 31, 112, -18, -83, 6, 125, 29, -83, 54, 111, -2, -83, -124, 25, -56, -102, -67, -20, -40, -64, -120, 9, -84, -64, 127, -4, -21, 54, -98, -42, -96, -126, -65, 78, -33, -88, -81, -62, -63, 58, 24, 66, -24, -94, -74, -15, -107, 72, 14, 66, 18, 17, 56, 35, 45, 96, 29, 20, -127, 40, -44, 48, 82, -51, -14, -108, -71, 126, 2, -38, 82, 28, 6, -27, 57, -39, 109, -30, 49, -84, 35, 87, 38, 106, -90, -99, 115, -67, 100, 0, 1, -66, 71, 63, -28, -57, 28, 6, -105, 88, 8, -61, 5, -27, -53, -112, 85, 68, 86, 122, 4, -81, -63, -50, -45, -74, 90, -78, -24, 46, 10, 72, 14, 29, 64, -101, -128, -73, 90, -16, -14, 13, 124, 12, 59, -96, -32, -10, -35, 116, 90, 61, -101, -56, 73, -96, 71, -41, -49, -39, 68, -126, -124, 59, -82, -73, 102, -12, -114, -14, 63, -15, -89, 121, 46, -112, 15, 78, -43, -60, 36, -67, 22, 106, -10, -49, 1, -14, 49, 46, -16, 35, -81, -4, -49, 41, 45, -92, -34, -54, -118, 52, -42, -9, 99, -14, -108, 57, 73, -14, 112, 122, 66, -128, 27, -90, 80, -26, -74, 30, 90, 48, 25, 64, -66, 75, 74, -85, 50, 60, 47, 106, 88, -124, 47, 101, -109, 4, 18, -11, 72, 91, -105, 112, -14, 121, 127, 75, -96, -65, -58, -11, -64, -40, 51, 93, -114, -1, 23, 18, -78, 46, -46, -37, 50, 28, -107, 57, 122, -54, 9, 7, 76, 11, 122, 58, -17, -114, 125, -10, 54, 8, 46, 84, -125, -124, -5, -56, -29, 11, -108, 14, 94, 103, -49, -39, 73, 74, -70, -83, -13, -12, 18, -89, 109, 97, -100, -34, 86, -80, 5, 12, 124, -64, 93, -72, 36, 123, 69, 41, -58, 82, -114, 43, 96, -123, -121, 21, 25, -100, 99, -53, 90, 119, -87, 15, 95, -84, -98, 11, -15, 108, -111, -15, 76, 84, 123, -116, 63, -24, 2, -121, -33, 78, 92, -109, 116, -65, -15, 9, 49, 85, -17, -28, -48, 97, -48, 70, -102, 8, -49, -101, -115, -32, 88, 80, -105, -4, 123, 26, -29, -54, -102, 89, 50, -13, 105, 84, -65, 53, 113, -106, -59, 9, -86, 95, 26, 74, -121, -70, 32, 45, 22, -106, -128, 80, -57, 41, -123, -11, -23, -125, -70, 50, -104, -12, -109, 30, -5, -20, -52, 62, -68, -88, 13, -98, -9, 6, 94, 97, 36, 110, -52, -19, 83, -7, -54, -45, 45, -23, -90, -98, -98, 79, 84, -67, 85, 2, -10, -78, 24, 56, -29, -40, -33, -40, -26, 48, 7, 101, -45, -41, 115, 24, -26, -63, 29, -58, 52, 58, 69, -36, -80, 75, -21, -93, -110, 89, -77, 48, -122, -25, -115, 7, -96, 91, -71, -23, -16, -59, 22, 121, -74, -89, -97, 49, -77, 33, -63, 39, 3, 59, 109, -59, 109, -94, 123, 4, -110, -127, -38, -11, 92, -18, 66, 67, 58, 56, 53, -107, 16, 107, -78, 52, -73, -94, 6, 34, -85, 76, -112, -94, -90, 58, -40, 37, -3, -77, -90, -102, -1, -79, 4, 38, 27, 111, -109, 8, 18, 120, -80, 3, 99, 5, -128, -62, 97, -27, 110, -111, 23, 74, 80, -92, -108, -17, -115, -83, 59, -3, -122, 37, -118, 54, -18, -88, 120, 67, -25, -87, 77, -35, -34, -14, -43, -58, 99, 115, 40, -85, -100, 79, 63, 115, 75, -48, 55, -20, 41, -75, -50, -27, -93, -2, -9, 35, 35, 75, -39, 109, -60, -73, -10, -62, -128, 90, -66, 13, -79, 74, -14, 108, -36, -89, -46, -45, 111, 0, -68, -14, -106, -5, -12, 52, 35, 10, 0, -1, 77, -14, -59, -54, -29, 34, 123, 116, 99, -32, -109, 15, -125, -78, 35, -119, -89, 81, 59, -116, -110, -70, 96, -22, -16, -38, 97, -35, 56, -61, -126, -103, -13, 85, 96, -7, 68, -113, -77, -105, -30, 0, -45, 69, 68, 32, 22, -117, 43, -46, 18, -94, 114, 37, 35, 94, 125, -52, -16, 15, 118, 25, -108, 118, -49, -126, -125, 27, -83, 95, 62, 2, -63, 95, 94, -54, -9, 82, 51, 28, -29, 46, 60, -4, 90, -86, -118, -74, 91, -63, 127, -104, -32, -2, 120, -69, -22, 28, 7, 101, -42, 95, 99, -127, 113, -89, -119, -89, 81, 50, -53, -3, 118, -35, 2, -23, 18, -19, -99, -96, 102, -114, 26, 75, -113, -4, 53, 95, -36, 18, -4, -64, -112, 49, 75, -73, -102, -58, 5, 64, -43, -25, -37, -1, -110, 44, 92, -85, -124, -128, 30, 3, 24, 71, 26, 107, -112, -37, 53, -113, 126, -35, 19, -53, -46, 83, -37, 70, 78, -109, -15, -85, -30, 3, 92, -92, -65, -109, -35, -96, 32, 105, 126, -13, 126, -89, -16, 74, -113, 23, -128, 85, 45, -11, -36, 9, -1, -38, 106, -109, -33, 80, -94, 85, 127, 56, -72, 116, -119, 76, 63, -123, -13, -103, 65, -2, -70, -70, 40, 87, 40, -103, 96, 23, -43, -69, -74, -30, -56, 125, 72, -42, 11, 71, -32, -6, 95, -40, -14, -12, -71, 119, 26, 13, 32, -80, -126, -58, -76, 107, -6, 15, 110, 13, 107, -36, -118, 36, 0, 89, 108, 53, 63, -68, -80, -38, 61, 59, -120, -6, 42, 39, 114, -38, 26, 85, 125, -120, -113, 101, -30, -43, -29, -65, -85, -41, 12, 9, -38, 100, -26, -29, -30, 95, -66, 88, 56, -61, -79, -78, -119, 124, -92, -10, 22, 67, 103, -27, 98, 9, 13, 87, -122, 59, 114, 6, -55, 59, 30, -5, 53, -76, -117, -86, -14, -13, -45, -92, 40, -16, -9, 52, 71, -65, 56, 97, -78, -100, 16, 39, -24, 117, -62, -126, -39, 108, 49, -88, -112, -13, -63, 56, 111, -45, -124, 96, 31, 14, -105, 23, -117, 11, 65, 23, 99, 27, -51, 73, 126, -44, 82, 23, -47, 17, -86, 92, 27, -27, -87, 47, -99, 21, 45, -8, -127, 88, 56, 102, 9, 83, -52, -104, -30, -9, 48, 116, -17, -69, -53, 75, -20, 86, 1, 80, -89, 56, 17, -81, -62, -99, 11, -7, 99, 108, -32, -21, -27, 92, 79, -98, 44, -61, -3, -106, 31, 57, 104, 88, -91, 36, -11, 79, 89, 126, -27, -124, 25, 9, -69, 125, -105, -29, 38, -99, -30, -60, 36, -52, 15, -104, 58, -122, -68, -101, 85, 25, 45, -128, 21, 30, 19, -81, -99, 34, -87, -79, -23, 58, 21, -108, 33, -124, -47, -46, 88, 96, -90, -28, 49, -116, 19, -56, -72, -43, -95, -120, -13, 6, -100, 26, 11, -72, 51, -100, -104, 64, 75, -21, -6, -127, -113, 9, -2, -92, -61, -24, -118, -91, -27, -53, -105, -69, 127, 109, 85, -126, 126, -66, -98, -83, 45, -44, 117, -120, 17, 108, -117, -7, -71, -78, 70, 48, -47, 74, 55, 69, -15, 0, 54, -92, 99, -109, 7, -9, 48, 106, -75, -26, 27, 26, 70, -63, -26, -75, 44, -81, -44, 0, -111, 83, 12, -116, 9, 58, -58, -14, -74, 8, -33, 0, 107, 65, 22, 84, -49, 36, -36, -12, -53, -40, -5, -114, 97, 84, 81, -2, 41, -41, -69, -110, 125, 31, -8, 57, -3, -96, 124, -12, -91, 7, -33, 15, -82, 20, 47, 10, -96, 67, 3, 3, -44, 77, 78, 63, -101, 2, 81, -5, 79, 21, -34, 79, -30, 106, 68, -95, 5, 120, 36, 24, 81, 5, 41, 74, -31, 117, -7, -23, -47, 114, 80, -8, -35, -122, 100, -8, -45, -79, 8, 96, 4, 105, -16, -94, 79, -36, 4, -53, 61, -99, -112, -69, 117, 69, 99, -7, 10, 13, 98, 60, 10, -2, 112, -112, -43, -79, 82, 47, 117, -116, 100, 77, 122, -57, -124, -63, 33, 42, 126, 58, -86, 97, -68, 61, -95, -79, -53, -27, -26, 48, 92, -42, 4, 98, -18, -110, -91, -64, -64, -10, -121, -50, -40, 104, 13, 75, -60, -107, -47, 95, -57, -58, -97, 66, 62, 116, -91, 125, -24, -112, -103, -17, 35, 80, -81);
    signal scenario_output2 : scenario_type2 :=(-57, -40, 46, 127, -40, -86, 26, -26, 115, -76, 8, 26, -64, 24, -94, 115, 121, -64, -119, 64, 76, -128, -68, 40, 72, -9, -10, -54, 70, 127, -128, -43, 103, -20, -128, 93, 74, -58, 89, -128, -88, 69, -55, 90, 72, -77, 22, 62, -37, -83, 54, -46, 17, 108, -128, 48, 116, 17, -68, 1, 108, -109, 26, 65, -114, -113, -25, 127, -46, -20, 104, -62, -49, 72, -10, -97, -15, 127, -18, -128, 127, 7, -122, -46, 127, 8, -128, 38, 119, 95, -128, -57, 127, 69, -111, 24, 48, -1, -104, -20, 23, -65, 127, -82, -66, 9, -9, 0, 78, 125, -128, -47, 14, -29, 93, 59, 27, -99, -122, 110, 32, 44, 30, -108, -49, 64, 104, 8, -77, -9, 0, 66, -41, -128, 7, 37, 127, -46, -61, 21, -40, 22, 2, 13, 113, -119, 21, -9, -37, 127, -82, -1, -70, 60, 24, -108, 123, -26, -3, -2, -12, 51, -115, -41, 3, -18, 53, 46, -8, -79, 14, 70, 97, -100, -128, 127, 96, -128, -83, 53, 14, 29, -28, 58, 0, -30, 62, -83, 35, -42, 86, 68, -128, 81, 76, -29, -36, 31, -30, -69, -2, 58, -82, -30, 12, -51, 99, -38, -55, 69, -9, -18, 82, 64, -94, -97, 127, -5, 8, 72, -128, -82, 127, 22, -128, 114, 100, -38, 71, -128, -48, 127, -97, -108, 77, 111, 12, -115, -116, 103, 122, -121, 3, 49, 5, -6, 6, 40, 5, -10, -111, 70, 72, -65, -42, 26, 110, -42, -128, 1, 126, 10, -42, -107, 45, 29, -24, 127, -128, -72, 127, -54, -58, 105, -123, -46, -2, 87, 11, -39, 127, -128, 11, 40, -128, 71, 39, 0, 22, 11, 49, 45, -64, -128, -10, 127, -88, 38, 52, -58, 113, -21, -55, -9, -48, 22, -45, 8, 127, -29, -128, -47, 4, 34, 24, -51, -44, 127, 85, -127, -62, 70, 127, 7, -128, 43, 77, -128, 4, 123, -73, 36, 115, -55, -128, 8, 127, 48, -57, -126, -29, 28, 40, -56, -40, 127, 8, -38, -13, 3, 31, 2, -64, -68, 38, 113, -14, 7, -27, 0, 38, 42, -44, -128, 72, 24, 15, 28, -19, 30, -35, -127, -39, 127, 8, -49, 42, -64, 91, -14, -11, 57, -86, 9, 43, -4, 55, -70, -53, 47, -13, -29, 37, -68, -104, 61, 70, 53, 62, -35, -37, 75, -96, 12, 18, -77, -40, 82, 89, -48, 24, 51, -110, -81, 127, -90, -107, 38, 73, 63, 38, 41, -128, -21, 112, -76, 59, -55, -35, 127, -126, 48, 106, -38, -36, 31, -45, -64, 19, -70, 11, 126, 51, -128, 104, -34, -128, 127, -42, -70, 98, -4, 53, -29, -128, -18, 127, 9, -128, 73, -24, 36, 127, -128, -128, 127, 25, -81, 21, -15, 54, -44, 1, 38, -19, -29, -11, 5, 13, 100, 42, -78, -109, 127, -55, 8, 18, -8, 68, -121, -46, -15, 127, 61, -128, 58, 127, -83, -105, -54, -46, 127, 57, -27, 28, -92, -9, 37, -40, 12, 17, 43, 26, 9, 23, -128, -5, 27, 95, -31, -66, 7, -55, 75, -59, 127, -26, -42, 42, -59, 7, -102, 89, 110, -57, 23, 12, -61, -83, 41, 127, -76, -98, 114, 98, -128, -128, 47, 115, 28, 0, -21, 21, -42, -128, 45, 63, 56, -66, -4, 81, 15, 36, -121, -109, 75, 127, -48, -128, 109, 127, -107, -93, -18, 51, 93, 18, -106, -73, 59, 28, 34, -42, -58, -12, 58, -1, -46, -3, 14, -10, -28, 6, 0, -3, 110, 13, 9, 85, -128, -44, 125, 31, 40, -128, -25, 127, 25, -62, -40, -61, -103, 87, 7, -80, 26, 98, -18, 11, 41, -81, 30, 114, -44, -71, -2, 19, -4, -10, 2, 40, -22, -128, 59, 52, -34, 91, -55, -41, 107, -69, -58, 81, 6, -120, 127, -36, -77, 127, -3, -29, -73, -64, 125, 93, -96, -73, -51, -30, 115, 13, -15, -20, 35, 28, -53, 100, -60, -89, 47, 32, 11, -14, 2, -98, 92, 8, -128, 88, 115, -47, 34, -18, -68, 55, -32, -46, 46, 39, 8, 72, -119, -94, 66, 5, 55, 85, -69, -127, 23, 122, -54, 19, 40, -128, 105, 90, -128, 57, -13, -71, 77, 13, -78, 52, 4, -70, 17, -27, 127, 64, -3, -74, -59, 127, -34, -127, 62, -37, -39, 36, 23, 13, 61, 0, -12, 20, -112, 12, 54, -100, 83, 106, -88, 40, -5, -79, 28, 30, -14, -66, 18, -1, -95, 42, 72, 15, -28, 22, -28, -51, 127, -15, -6, 104, -27, -108, 24, -28, 36, 74, -71, 2, 46, -1, 4, -30, -79, 82, -7, 14, 59, -30, -46, -117, 63, 120, 17, -109, -128, 58, 63, 112, -94, -29, 127, -128, -119, 110, 113, -82, -5, 127, -128, -99, 60, 46, 6, -94, -29, 35, -31, 17, 105, -57, -36, 5, -42, 27, 45, 66, -111, 23, 38, -87, -14, 105, 112, -83, 68, -89, -102, 127, -96, -81, 98, 21, -2, -99, 98, 10, -41, -9, -128, 127, 70, -103, 14, 94, 21, -128, -6, -24, -10, 9, -6, 77, -22, 85, 52, -42, -128, -9, 122, -102, -34, 127, -13, -91, 59, -18, 66, -56, 8, -27, -24, 80, -95, 83, -57, -112, 127, 127, -75, -105, -18, 4, 8, -54, 38, 70, -37, 94, -14, -22, 54, 24, -61, -55, 63, 22, -100, 28, 115, -68, -91, -3, 56, 0, 18, 12, 73, -128, -54, 94, -76, 5, 14, 10, -42, 43, 24, -116, 2, 127, -78, -28, 127, -5, -18, -20, -12, -123, 81, 42, -128, 23, 120, 34, -76, 37, -44, 47, 29, -75, -15, -30, 69, 24, -42, -40, -26, 62, 52, -114, 94, 76, -126, 41, 4, -61, -39, 49, 8, 1, 98, -128, 3, 89, -62, -66, 112, 44, -24, 106, -128, -74, 11, 71, 15, -78, 32, 34, -32, 52, -44, -126, 127, 52, -66, -85, 127, -3, -128, 105, 97, -90, 19, 13, 30, -17, -54, 44, -37, 56, -49, 0, 113, -107, 22, 111, -128, 19, -18, 31, 127, -128, 25, -23, -97, 127, -59, -31, 92, -20, -31, 70, -22, -34, 74, -29, -104, -23, 127, -76, -11, 127, -59, -60, 95, 71, -55, -2, -92, -93, 56, 109, 99, -128, -52, 116, -112, 106, -39, -28, 127, -90, -62, 80, 19, -124, -69, 83, 30, -17, 62, -38, 0, 2, 2, -53, 40, 5, -43, -30, 18, 127, -52, -128, 55, 127, 17, -60, -64, -24, -35, 98, 9, -63, -75, 56, -9, -32, 127, -43, -120, 127, -34, -27, 123, -6, -115, -87, 59, -28, 6, 46, 90, -53, -112, 112, 72, -128, -58, 6, 52, 126, -19, 32, -36, 27, -53, -63, 9, -109, 66, 110, -14, -80, 113, -28, -19, -40, 34, 91, -46, -95, 41, 127, -128, -60, 24, -34, -58, 93, 42, -32, 70, -119, 79, 52, -85, 15, -77, 43, -17, 65, 4, -82, 29, -43, 41, 1, 100, -15, -98, 38, -15, 29, 95, -28, -24, 14, -108, 11, -35, 57, 44, -76, -8, 56, -57, 72, 81, -42, 29, -95, -76, 127, -15, -38, 46, -8, 12, -103, 22, -19, 93, -20, -46, 25, 4, 60, 30, 8, -128, 54, 127, -71, -19, -5, -61, -56, -5, 32, 9, 89, 109, -105, -128, 127, 48, -128, 64, 123, -122, -58, 114, -78, -12, 76, 21, 9, -10, 46, -85, -31, 59, 38, -19, -128, 64, 17, 38, 103, -44, -128, 107, 13, -128, 60, 30, -45, 106, -22, -19, 127, -20, -104, -128, 127, 65, -128, -31, 127, 29, -77, -66, 97, -64, -5, 127, -1, -72, -19, 127, -128, -1, 127, -65, -128, -71, 83, 17, -89, 78, 69, 73, -98, -44, 107, 20, -128, 44, 65, -128, 47, -39, -31, 75, 75, -96, 70, -10, -66, 127, -51, -99, 116, -28, -128, 127, 11, -2, -1, -128, 123, 26, 27, -49, -45, 61, -25, -7, -11, 121, 15, -7, -49, -8, -97, 29, 127, -70, -53, -2, -80, -60, 45, -15, -40, 29, 6, 100, 87, -128, 2, 44, -74, -37, -12, 110, 34, -111, -57, 110, 100, 6, -63, -64, -26, 29, 6, -60, 45, 35, -32, 105, 31, -120, 28, 37, 61, -45, -47, 97, -30, -47, 26, -44, 57, -29, -124, -8, 48, -10, -34, 104, -23, 35, 47, -10, 14, -55, -70, -70, 100, 30, 61, 12, -111, 78, 46, -30, -32, 4, -34, 83, -89, -3, 127, -128, -11, 106, -97, -5, -1, -53, 75, 45, -119, 105, 14, -128, 93, -34, 51, -6, -49, 26, 86, -32, -95, 127, -89, -105, 12, 80, 106, -128, 42, 114, -128, 78, 127, -128, -3, 61, -37, 94, -96, -45, 102, -63, 49, -28, -128, 22, 45, 7, -6, 14, 8, -110, 97, 127, -17, -128, -7, 127, -36, -52, -25, 39, -83, 43, 113, -90, 18, -27, 68, -8, -21, 73, -128, 15, 120, -128, 38, 127, -128, 9, 35, -71, 20, 35, 51, 18, -43, -107, 127, 26, -94, 98, -71, -128, 127, -11, -6, 127, -128, -8, -4, -29, -15, 81, 34, -128, 59, 61, -62, -71, 100, -1, -54, 1, 63, 127, -89, -42, 77, -93, 8, 1, -52, 127, -42, -32, 3, -65, 89, 53, 34, -120, 36, 19, -128, 32, 97, 20, -57, -32, 4, 94, 1, -117, -69, 60, 6, -61, 127, 47, -103, 111, 26, -128, 80, 74, -36, -83, -25, 86, 22, -64, -94, 47, -31, 112, 13, -128, 126, 123, -113, -125, 127, 45, 36, -88, -34, 127, -62, -121, -98, 77, 122, -38, 2, -10, -51, 90, 22, -89, 72, -10, -106, -41, 61, 111, -122, -47, -21, 126, 14, -128, 127, -13, -5, 11, 0, -22, -81, 122, -34, -59, 127, -70, -6, 23, -128, 104, 127, -128, 5, 53, -57, 25, 48, 41, -113, -17, 116, -20, -38, 48, -61, -26, 42, -121, 87, 29, -27, 124, -35, -1, -99, -5, 28, -56, -6, 74, 76, -46, 96, -128, -22, 73, 19, -57, -100, 69, 55, 106, -128, -36, 17, 6, 127, -59, -30, -74, -30, 127, -1, 19, -8, -128, 26, -20, -71, 65, 112, 83, -53, -128, 0, 127, -35, 13, 73, -92, -126, 83, 127, -42, -99, 28, -45, -96, 34, 0, 61, -17, -40, 127, -3, -127, 23, 37, -30, -31, 77, -5, -96, 28, 41, 107, -62, 3, -32, -65, 60, -106, 96, 2, -80, 42, -11, -19, 32, 74, 9, 55, -26, -128, 79, 22, -114, 127, -29, -1, 51, 4, -54, -47, 62, -21, 68, 17, -79, -24, -34, -66, 41, -31, 94, 57, -23, -86, 21, 127, -1, 9, -45, 24, -90, -123, 127, -49, -28, 51, -109, -47, 127, 66, -29, 86, -82, -95, -34, 127, -4, -128, 64, 36, 64, -77, -39, 36, 70, -41, -98, 109, -43, -61, -11, 103, 79, -49, -105, 46, 96, -22, 59, -30, -106, -29, 29, 48, 48, 60, -127, -14, 19, -22, -9, -55, 6, -29, 94, 127, -64, -114, 127, -11, -51, -5, -77, 0, 0, -27, 63, 127, -25, -21, 11, -34, -60, 12, 127, -107, -37, 116, -37, -7, -103, 49, 0, 39, 0, -75, 41, -81, 108, 40, -38, 0, -68, 115, -69, -119, 96, 66, -102, 47, 4, -1, 45, -79, 127, -120, 0, 127, -128, -95, 73, 41, -4, -37, 44, 17, -62, 27, 40, 8, 0, -6, -73, 48, 91, -19, -115, 32, 23, -21, -68, -24, 79, -89, 62, 83, -30, 45, -108, -85, 127, 43, -87, 36, 11, -81, -35, 75, -40, -78, 81, -27, -47, -44, 127, 127, -73, 3, -52, -128, 27, 82, 72, -36, -4, 77, -28, -105, 66, 43, -49, 37, -15, -9, -66, -34, -20, 9, 44, -38, 64, -46, 4, 81, -38, 2, 65, -86, -6, 76, -128, 66, 3, -54, 8, 106, 41, -108, 20, 93, -28, -99, -13, -18, 92, 88, -103, -34, 39, 31, -56, 1, 127, -128, -47, 60, 54, -20, -128, 127, 119, -128, 60, 107, -128, 28, -25, 32, 26, -44, -2, -19, 93, -115, 9, 46, -35, 60, -52, 18, 117, -109, -95, 127, 46, -115, 11, -29, -15, -18, 60, -2, 43, -21, -63, 60, -37, 1, 74, -24, -5, 35, 12, -87, 8, 44, -74, 127, -40, -128, 53, 68, -29, -14, -49, 17, -18, -35, 47, 0, -70, 102, 123, -2, -98, -114, -7, 105, 55, -74, 79, 107, -64, -94, -36, 41, 127, -127, -49, 86, -8, 14, -80, 89, -7, -49, 121, -56, 36, -91, -4, 63, -78, 73, -26, 21, 23, -106, 76, 11, -43, 103, 34, -102, -108, 66, 121, -110, -100, 43, 74, -20, -72, 57, -42, 20, 104, 15, -56, -21, -83, 9, 127, -95, -56, 93, -123, 72, 47, -2, -44, 28, 18, -53, -6, -73, 109, -29, 66, 4, -128, 94, 20, -124, -25, 8, 127, 37, -73, 57, 56, -99, -93, 7, 91, 99, 12, -110, -66, 18, -30, 10, 97, -6, 29, 14, -32, -5, 29, -3, -110, 18, 98, 94, -100, 0, -45, -30, 97, -61, 46, -65, -43, 127, -127, -10, 80, -108, 32, -62, 62, 98, -65, -7, 13, 74, -46, -32, 102, -10, -126, 8, 127, -107, -128, 12, 24, 127, 0, -24, -10, -66, 125, -52, 8, -3, -119, 2, 41, 90, 4, 52, -128, 29, 127, -78, -122, 79, 63, -85, 77, 56, -36, -25, 31, -105, -38, 30, -43, 69, -54, -119, 127, 96, -74, -36, 75, -55, 18, 125, -85, -54, -92, 44, 100, 12, -30, -102, 71, 81, 1, 0, -128, 41, 127, -128, -95, 44, -31, 27, 120, -4, -66, 72, 45, -79, 47, -26, -56, 19, -87, 92, 125, -120, -99, -23, 98, 122, -29, 5, -27, -5, -55, -104, 105, -36, -62, 117, -37, -26, -14, -37, 105, 7, 37, 77, -5, 11, -128, 38, 18, -65, 127, 13, -22, 7, 81, -128, -103, 127, -24, -128, 64, -5, 34, 81, -128, 86, 15, -103, 127, 3, -87, 28, -40, -88, 49, 127, 0, -128, -63, 83, 68, -37, 54, 51, -126, -44, 92, -60, -61, -35, 104, 58, -116, 92, 96, -5, 12, -87, -49, -29, -74, 110, 104, -27, -128, -6, 95, 66, -56, -128, 45, 127, -97, -95, 37, -77, 28, 112, 4, -120, 83, 52, -123, 13, 127, -83, -100, 127, -45, -62, -18, -44, 85, -9, 34, 116, -39, -128, 105, -17, -98, 52, 54, 119, -80, -100, 108, 18, -29, 76, -110, -4, -13, -128, 109, 127, -90, 3, -43, 41, 85, -72, -21, -6, 104, -113, -83, 19, 112, 15, -128, 127, -21, 2, 25, -128, 107, 88, -73, 64, -73, 0, 96, -57, -76, -69, 114, 51, 3, -83, 39, 35, -128, 105, -36, -21, 127, -97, 64, -4, -128, 127, -55, -127, 127, 104, -128, -8, -32, 25, 113, -128, -1, -10, 93, 98, -126, 10, -4, -13, 7, 27, 0, -112, 70, 106, -25, -128, 56, 44, -27, 25, -54, 7, 28, -62, -88, 127, 76, -6, -70, 1, 23, -128, 7, 79, -6, -45, -19, 81, 127, -99, -25, -10, -2, -37, 34, 35, -60, 92, -61, -3, 58, -94, 24, -1, -13, 80, -66, -38, 41, -65, 59, -18, 43, 21, -43, 7, 23, 127, -114, -74, 62, -72, -49, 9, 105, 127, -61, -128, 18, 94, -15, -98, 72, -11, -80, 127, 52, -128, -29, 103, -12, 41, -128, 46, 127, -128, -55, 57, -80, 87, 127, -128, -128, 127, -7, -19, 127, -128, -115, 111, 11, -37, 55, 40, -24, -76, 6, 114, -73, 25, 61, -7, -39, 19, -40, -70, 110, -15, -7, -12, -72, 26, 127, -128, -30, 96, -128, 74, 90, -44, -63, 14, 49, -30, 18, -82, -8, 127, 0, -127, -79, 53, 38, -82, 82, -23, -5, 54, -35, 107, -46, -128, 127, 81, -97, 54, 22, -119, -40, 127, -30, -52, 15, 47, -13, -128, 9, -20, 124, 6, -38, 75, -105, 35, 55, -23, 0, -43, 10, 61, 41, -128, 47, 26, -43, 127, -17, -92, -19, -6, -112, 97, 127, -9, -122, -69, 59, -46, 83, -26, -82, 47, 49, 100, 0, -11, 15, -89, -122, -4, 127, -27, -54, 127, -77, -60, 127, -81, -128, 127, 39, -27, -44, -59, -18, -29, 0, 127, 34, -81, 46, -124, 53, 83, -34, 14, -95, -56, 127, -48, -107, 122, 34, 6, 51, -121, 24, 78, -28, -80, 14, 108, -128, -106, 127, 25, -128, 127, 29, -90, 45, -49, -47, 46, -20, 30, -37, 56, 127, -94, 44, -20, -120, 49, 114, -85, -91, 91, 43, 36, -17, -19, -77, 43, 77, -52, 77, -128, 5, 113, -100, -75, 28, 9, -36, 18, 48, -63, 43, 60, -2, 11, -73, 21, 80, -49, -25, 127, -128, -23, 94, -86, -51, 112, -11, -128, 127, 4, -23, 109, -44, -63, -120, 31, 86, -42, 51, 13, -25, 63, -70, 36, 94, -42, 11, -54, -115, 74, 127, -41, -97, -62, 69, 87, -47, 37, 57, -128, 45, 34, -128, 127, 127, -29, -128, 15, 127, -128, 40, -36, -30, 36, -128, 127, 112, -51, 26, -79, -79, 122, -70, -109, 127, 40, -11, -93, -58, 91, 14, -106, 12, 95, -111, 0, -17, -21, 127, -46, 0, -19, -78, 127, -42, -57, -54, 26, 82, -14, 8, -10, 9, 70, 32, -97, -22, -6, 14, -38, -5, -39, 55, 78, 21, -35, -110, 79, 3, 66, -55, -21, -46, -5, 115, -39, 11, -92, -82, 39, 22, 2, -32, 53, 102, -65, 47, -64, -38, 68, -18, 92, -24, -65, -36, 56, 31, -47, -59, -18, -7, 111, 87, -41, -26, 22, -1, -117, 108, -39, -128, 53, -17, 70, 6, -112, 107, 19, 69, -15, -77, 61, 31, -94, -32, 127, -128, 68, 20, 6, 28, -60, 127, -119, -81, 74, -58, 19, 45, 65, 19, -128, 48, 4, 19, 36, -53, -26, 57, 0, -51, 116, -128, 22, 127, -128, -68, 12, 80, 93, 3, -126, -68, 43, -57, 31, 46, 59, -63, 20, 127, -111, -79, 34, -56, -17, 3, 70, 120, -80, -29, -8, -20, 127, -35, -104, 10, 99, -63, -110, 6, 35, 75, -52, -14, -15, 40, 57, -88, -9, -18, 102, 49, -10, 43, -10, -11, -97, 56, 64, -128, -18, -44, 124, 5, -128, 127, 86, -5, -45, 13, -106, 21, 68, -128, 113, -18, -8, 90, -10, 0, -128, -11, 52, 46, 56, -128, -52, 26, -23, 10, -25, 100, 117, -43, -94, 92, 9, -128, 21, 42, 27, 82, -45, -128, 79, 60, -34, -24, 22, -7, -51, 4, 19, 40, 14, -65, -21, 116, 9, -40, 52, 27, -53, -39, -47, -5, 68, 88, -36, -117, 30, -3, -40, 113, 47, -99, -98, 35, 91, -61, -34, 127, -6, -128, 17, 127, -108, 42, 31, -32, -38, 2, 127, -79, 34, -113, -1, 39, -51, 85, 35, -12, -128, 106, 22, -89, 127, -90, -128, 55, -11, -2, 68, 56, -69, 19, 28, 14, 71, -128, 22, 109, -54, -89, -54, 127, 40, -117, 53, 6, -74, 127, 127, -124, 5, 72, -52, -76, -78, 83, 112, -41, 4, -102, 3, 64, -24, 34, 37, -104, 8, 41, -95, 71, -2, -34, -86, 127, 25, -36, -3, -94, 46, 79, -51, -116, 24, 89, 111, -99, -38, 117, 8, -42, -58, -24, -61, 61, -13, 28, 127, -128, 52, -11, -119, 106, 108, -37, -39, 56, -111, 7, -8, -19, 125, -97, -1, 58, -97, 1, 1, 15, -22, 2, 79, -64, -14, 109, -79, -60, 93, 122, -113, -1, 94, -92, 44, 52, 2, -23, -70, -68, 48, 0, -48, 23, 64, -55, 29, -5, -29, 127, -107, 14, 127, -38, -128, -59, 93, 71, -22, 13, -59, -44, 115, -102, -103, 90, 32, -71, -11, 31, -30, 99, -19, -105, 28, -25, 49, 127, 19, -128, 61, 83, -128, 109, 97, -66, 55, -88, -21, 115, -81, -58, 24, -51, 105, -49, -73, 25, -41, 72, 64, -58, 13, 88, -110, 47, -25, -8, -24, 61, 14, -64, 77, -52, -8, -73, -28, 77, 74, -47, -113, 127, 30, -128, 127, -51, -69, -11, 2, 65, 53, -69, -27, 63, -69, 1, 23, -42, 47, 27, -112, 11, 62, -17, -88, 116, 121, -69, -19, -46, -60, 65, 9, -31, -3, -63, 99, 127, -128, 31, -29, -30, 59, -128, 103, 69, -103, 85, 5, -116, 4, 0, 77, 82, 42, -14, -128, -73, 83, 29, -73, 31, 110, -34, -128, 55, 68, -54, -13, 48, 69, 14, -42, -42, -66, 31, 93, 11, -119, 39, -20, -7, 82, -128, 124, 0, -27, 127, -103, -62, 25, -88, 14, 127, -49, -4, 99, -45, -75, 70, 19, -19, -2, -96, 1, 122, -96, -29, 127, -8, -52, 24, -68, 18, 127, -128, -19, 111, -107, 25, 127, -128, -94, -11, 71, 96, -128, -58, 107, 12, 77, -65, -126, 104, -3, -89, 99, 62, 41, -91, -93, 127, -17, -128, 38, -14, -96, 127, -14, -109, 102, -61, 35, 0, -60, 82, -73, -55, 56, 86, 43, -107, -65, 53, -13, -48, 127, 4, -1, 27, -128, 127, 11, -128, 34, -39, 14, 62, -2, -81, 42, 66, 64, -43, -128, 127, 32, -34, 92, 0, -95, 37, 14, -76, 21, -64, -51, 63, -27, 74, 61, -20, 71, -43, -53, -86, 31, 20, 82, 73, -128, -36, -25, 10, 81, 34, -78, 51, 75, -60, 19, 62, -82, 13, 22, -128, 61, 64, 24, 14, -29, -25, 55, -47, -128, 127, -30, -57, 120, -47, 66, -39, -128, 77, 59, -2, -35, -107, 116, 112, -115, -95, 108, 17, 6, 20, -65, -11, 68, -45, -38, 91, -35, 42, 52, -58, 19, -18, -55, 13, -76, -20, 96, 75, 22, -52, -128, 127, -32, -128, 23, 47, 14, -81, 38, 55, -19, -32, 105, 49, -60, 48, -119, 17, 127, -108, -86, -6, 81, 19, 56, 82, -34, -92, -45, -25, 1, 85, -17, -77, 45, -48, 56, 113, -79, -26, 15, -10, -31, 17, -10, -39, 64, 62, 32, -1, -99, -52, 91, 47, -124, -95, 127, 127, -128, -110, 55, 8, -21, -42, 57, 54, -89, 46, 58, -79, 100, 89, -44, 20, -8, -1, -122, -66, 23, 25, 44, 85, 8, -15, 79, -94, -128, 123, 6, -110, 17, 19, 25, -88, 19, 127, -46, -62, 104, 34, -17, 22, -5, -116, 13, 110, -68, 31, 27, -82, -28, -77, 28, -24, 107, 35, -128, -26, 127, 30, -106, 70, 47, 9, -38, -55, 44, 92, 24, -31, -23, 46, -97, -41, 59, -17, -94, 70, 10, -80, 77, 18, -112, 58, 127, -128, 32, 86, -79, -47, -32, 19, -32, 127, -32, 32, 5, -107, 124, 66, -128, 19, 60, -61, 107, 29, -15, -20, -71, -72, -30, 34, -35, 74, 98, -128, 36, 100, -87, -17, 116, 62, -128, -8, -20, -35, 127, -39, -42, 105, -91, 5, 127, -79, -128, -47, 122, 12, -89, 15, -9, -4, 47, 43, -89, 26, 53, -2, -29, 18, 91, 5, -126, 14, 127, -72, 12, -55, -126, 127, 36, 1, -63, -92, 9, 63, 127, -128, -87, 82, -95, 92, 58, 5, -59, -6, 115, 30, -128, -8, 127, -56, -62, 13, 19, 57, -75, -128, 83, 60, -46, 63, 5, 1, 0, -7, 8, 0, -61, -80, 125, -70, -10, 73, 18, 36, -51, -2, -34, 47, 60, -43, 27, 8, 11, -114, -64, 88, 66, -128, 49, 12, -13, 2, -90, 98, -21, -18, -70, 55, 127, -4, -80, -56, 29, 24, -29, 70, 43, -128, 68, 4, -62, 42, -20, 64, -113, 18, 127, -71, -28, -22, 34, 51, -128, 59, 43, -9, 123, -102, 12, 66, -128, -100, 114, 7, -34, 109, -71, 42, 109, 3, -65, -32, 56, -95, -23, 98, 37, -93, -128, 58, 24, -24, 66, -38, 46, 36, -73, 1, 31, 34, -110, 89, 54, -128, 95, 40, 15, 0, -90, -2, 42, -66, 46, 46, -45, -18, 75, -25, -37, 127, -77, -85, 1, -35, -55, 24, 87, 45, -10, -104, 77, 86, -37, 44, -26, -106, -35, 120, 63, -72, -72, 106, -14, 4, -34, -125, 127, 77, -128, 34, 44, -128, 32, 94, 103, 0, -128, -68, 46, 51, -49, 10, 127, -24, -42, 48, 22, -57, -109, 10, -27, -13, 90, -72, 18, -23, 80, 15, -68, 110, -57, 56, -5, -128, 127, 3, -36, 115, -58, -40, -54, -74, 41, 81, -38, 48, -65, -10, 23, -9, 103, -42, -105, 10, 105, 65, -25, -94, 1, 76, -88, -23, 127, -27, -79, 30, -73, -3, -3, -31, 127, 41, -25, -100, 4, 59, -49, -41, 15, 5, -14, 66, 27, -38, 40, 106, -128, -27, 99, -55, -100, -26, 127, -29, 9, 9, -128, 44, -3, 98, 36, 0, -44, -37, 99, 7, -15, -76, 104, -27, -93, 36, 65, -36, -23, 123, -127, 7, 42, -94, 46, 30, -66, 62, 40, -62, 93, -103, -97, 73, 59, -12, -53, 113, -49, -128, 126, 127, -128, -64, 85, -55, -57, 102, 81, -116, -69, 76, -51, -83, 127, -2, -128, 62, 4, -61, 127, -7, -128, 127, 43, -128, -6, 127, -30, 1, -2, -128, -26, 47, 27, 75, 66, -7, 9, -124, 69, -18, -79, 24, -58, 21, 76, -79, 69, 81, -36, 64, -128, -22, 127, -31, 18, -53, -43, 76, -45, 57, -7, -81, -82, 39, 28, -19, 127, -21, -20, 3, -15, 42, -128, -26, 53, -59, 17, 6, 88, 92, -128, -114, 94, 86, 23, 15, 6, 26, -81, -77, -72, 70, 112, -72, 8, 10, 45, -53, -65, 127, -93, -53, 127, -5, -128, -56, 48, 61, 27, 35, -64, -91, 73, 36, -6, -78, -57, 102, 127, -105, -75, 65, -36, -9, -6, 105, 10, -83, 106, -29, -96, -52, -15, 57, 8, 85, 51, -10, -32, -92, -37, -34, 103, 127, -106, -55, -62, 44, 56, -53, -47, -1, 127, 46, -128, -32, 127, -11, -95, -96, 127, -6, -15, 22, -9, 88, -128, 70, 4, -12, 72, -111, -31, 82, -56, 41, 93, -91, -73, -51, -15, 72, 10, -20, 38, -66, 7, 64, -53, 104, 89, -38, -22, 8, -85, -64, -5, 59, 9, -128, 126, 69, -45, 82, -81, -65, 119, 94, -128, -54, 127, 19, -88, -76, 43, -69, 65, -9, -128, 127, 107, -128, 44, -28, -85, 127, 4, -128, -6, 65, 2, -35, -56, 30, 112, 6, -37, 24, -60, -15, 12, -53, -19, 90, 1, -42, 125, -4, -37, 44, -128, -26, 124, 53, -35, -49, 25, -93, -44, 57, -4, 32, 5, 6, 12, -56, -22, 62, -5, -41, 94, -11, -21, 24, -19, -15, -82, 0, 57, 89, -63, -1, 36, -25, 115, -72, -60, -26, -85, 12, 127, 31, -35, -9, -48, 92, -59, -117, 127, -37, 36, 55, -25, -88, 35, 98, -124, 98, -11, -76, 117, -55, -111, 55, -71, 36, 127, 38, -106, -44, 127, -72, 9, -70, 30, 64, -46, -59, -105, 127, 127, -128, -45, 127, -24, 1, 15, -82, -9, 70, 28, 7, -83, 39, 90, -128, -69, 52, 105, -85, -77, 57, -111, 127, 127, -90, -94, 71, -47, 9, 127, -128, 0, -48, -24, 13, -86, 102, 32, 24, 88, -91, -128, 25, 127, -36, -127, 55, 69, -21, -54, 7, -8, -56, 81, 70, -79, -66, -2, 62, -19, 30, 58, -32, 9, 12, -39, 27, -45, -72, 81, 120, -22, -115, 24, 40, -99, -85, 97, 127, -128, 8, 62, -128, -32, 78, -6, 25, 127, -128, -128, 127, 29, -61, -13, 0, 125, -86, -47, 127, -47, -128, 113, 127, -8, -109, -22, 83, -128, 21, 3, -104, 114, 76, 28, 26, 1, -128, 4, 85, -20, -46, -54, 2, 0, 15, -5, 74, -51, -75, 88, 95, 10, -82, -112, -4, 127, -71, 5, 100, -128, 36, -9, -48, 127, -75, -12, -18, 20, 0, 15, 32, -74, -12, -4, 36, -1, 127, -69, -22, -32, 8, 98, -123, -75, 36, 37, 6, -59, -28, 85, 35, 24, -4, -6, 38, -68, 32, -42, 41, -2, -96, 10, -20, 11, 30, 19, 35, 100, -89, -111, 28, -22, 31, -17, -48, 81, 100, -91, -128, 79, 127, -54, -122, 1, 96, 127, -128, 5, 127, -114, -57, 124, -64, -15, 127, -128, -66, 17, 117, -11, -128, 46, 11, 12, 9, 127, -56, -128, 127, 127, -106, -109, 112, 71, -38, -42, -99, 25, 13, -104, 127, 104, -81, 51, 54, -128, 0, 51, -47, 78, -3, -70, -21, 87, -66, -128, 127, 79, -9, -90, -41, 114, -25, -81, 37, 113, -97, 35, 69, -89, 98, -68, -4, 25, -110, 49, 77, -37, -55, 3, -40, -35, 65, 0, -54, 0, 94, 27, -31, 43, -77, 36, 79, -38, 17, -55, -42, -23, 9, 65, -30, 74, -3, -29, -29, 18, -35, -42, 127, -81, 12, 15, -12, 95, -77, -5, -74, 2, -12, 42, 21, -82, 105, -27, 0, 68, -91, 2, 0, -102, 127, -32, 7, 72, -47, 9, -59, -61, 4, -5, 41, 52, 2, -44, -26, -5, -1, 48, 111, -69, -72, 19, -26, -19, 30, 122, -112, -69, 127, -80, 58, 26, -91, 127, -104, -108, 63, 83, -11, -115, 69, 115, -19, -9, -44, -125, 100, 127, -43, -65, -28, 40, 14, -1, -117, -22, 127, 22, -128, 93, 13, -2, 37, -128, 105, -48, 20, -13, -121, 127, 12, -11, -14, -9, 54, 0, -82, -11, 19, 15, -3, 4, 107, -27, -68, 70, -26, -57, 90, -32, 2, 63, -43, -81, -40, 56, 105, 9, -125, -71, 38, 127, -23, -128, 17, 3, -49, 127, 89, -119, -63, 110, 100, 18, -128, -63, 23, -83, -7, 127, 34, -44, 21, -22, 58, 76, -110, -103, 52, 113, -111, 30, -7, -68, 39, 49, -17, -128, 127, 71, -128, 38, 127, -97, -107, -4, 58, -18, -49, 28, 37, 40, 40, 34, -80, -5, 75, -92, 0, 103, -43, -79, 2, -51, 107, -19, -77, 96, -78, -76, 125, 127, -90, -34, -18, -52, 127, -65, -128, 71, 127, -85, -63, 127, 15, 17, -115, -34, -40, 75, 97, -128, 85, 94, -122, 23, 10, 41, 48, -110, 0, -79, 79, 63, -128, 72, -24, 23, 127, -128, 1, 127, -113, -29, -18, 0, 127, 48, -127, -108, 123, -73, -2, 127, -107, -105, 120, 39, -107, 64, -3, -88, 43, -62, -75, 82, -6, -37, 127, -10, -128, -35, 127, 36, 52, -77, -72, 79, -2, -56, -51, 127, -70, 8, 57, -86, -51, 0, 127, -88, -103, 127, 42, -52, -32, -35, 35, -39, 73, -35, -102, 5, 105, 114, -128, 36, 127, -34, -54, -89, 36, 79, -22, -112, 30, 127, -128, 36, 70, -46, 88, -128, 30, 127, -128, -6, 52, 39, 27, -128, 28, 127, -61, -111, 121, 106, -128, -5, -19, -52, 121, 76, -117, -81, 127, -27, -29, 25, -75, -53, 88, -18, -6, 30, -126, 111, 127, -96, -128, 27, 127, 48, -86, 22, -27, -46, -15, 35, 110, 12, -111, 18, 127, -56, -26, -54, 75, -76, -115, 92, -53, -49, 108, 55, -41, -36, -36, 52, 35, -85, 22, -11, 80, 0, -128, -3, 114, 127, -123, -62, 71, 77, -60, -128, 43, 103, 52, -45, 21, -41, -63, 124, 1, -93, -90, 65, 89, -43, -19, -35, -85, 53, 127, -83, 27, 26, -78, 127, -63, -108, 48, 98, 21, -128, 36, -26, 14, 110, -43, -70, -89, 83, -41, 112, -32, -40, 48, -112, 0, 81, 11, -83, 83, 56, -92, -6, 30, 79, 9, -128, 1, 28, -58, 127, 68, -128, 82, 104, -127, -2, 64, -128, 76, 127, -128, -57, -1, 72, -32, -65, 127, -87, -43, 51, 41, 28, -128, 55, 13, -83, 105, -31, 19, 89, 32, -56, -55, 93, -82, 8, -26, -72, 105, -37, -3, -63, 18, 127, -49, -85, 51, 4, -22, 48, 7, -119, 58, -11, 42, 2, -128, 127, 13, -20, 127, -121, -92, 72, 2, 91, 6, -128, 116, -43, -65, 98, 24, 32, -128, 64, 35, 25, -54, -88, 119, -64, 3, 48, -35, 1, 58, -71, 32, 94, -123, -78, 110, 15, -105, -57, 127, 68, -38, -54, -71, 127, -55, -106, 63, -57, 54, 10, 21, 104, -128, -106, -15, 127, 103, -62, -20, -81, -58, 100, 6, -34, 11, -44, -22, 97, -27, -95, 127, 47, -15, -52, -54, 127, -40, 8, -31, -117, 14, 85, -20, -71, 127, -55, -19, 46, 14, 93, -61, -97, -8, 30, 73, 76, -49, -29, 85, -96, -68, -15, 11, 74, -36, -59, 30, -34, -68, 127, -60, -113, 15, 105, 45, -42, 87, -79, -17, -58, 34, 10, 10, 14, -128, 126, -34, -49, 126, 31, -59, -1, 47, 1, 22, -30, -112, 44, -55, 47, 97, -125, 60, 0, 39, 14, -89, -27, 68, -72, -27, 21, 28, 3, 27, -7, -79, 68, -100, 82, 24, -86, 127, -21, -128, 127, -9, -57, 112, -115, 34, 120, -26, -76, -37, 27, 88, 6, -75, -62, -38, 88, 111, 5, -128, -45, 76, 53, -54, 1, 38, 13, 64, -128, -73, 114, -4, -106, 102, 82, -1, -100, 41, -29, -47, 112, -128, 5, 64, 3, -55, 97, 45, -45, 4, -51, 90, -44, -115, -19, -22, 85, 31, 74, -56, -28, 31, 0, -28, -107, 44, -10, 12, 123, 94, -128, 46, 18, -87, 73, -62, -32, 35, 75, -78, 60, 42, -128, 8, 46, -19, 61, -42, 30, -31, -18, 1, -13, 127, -73, -17, -13, 62, 10, -125, 20, -30, 79, 113, -90, -22, -37, -79, 90, 82, -61, 22, -53, 45, 127, -128, -41, 115, -27, -21, 7, -62, -48, 120, -21, -43, 80, -123, 59, 61, -128, 115, 24, -128, 44, 109, 25, -5, 59, -128, -47, 23, -86, 114, 68, -58, 85, -59, -48, 72, -12, -1, 36, -59, -107, 3, 77, 44, -72, 72, -45, 12, 127, -128, 11, 22, -107, 127, 120, -128, -119, 56, 7, 8, 52, 41, -10, -116, 38, 25, 68, 104, -128, 54, 36, -90, 69, 9, 85, -88, -109, -39, 96, 29, -102, 30, 70, -59, -30, 35, 82, 127, -128, -102, 127, -65, 14, 127, -128, -35, 21, -69, 112, -38, 38, 115, -62, -121, 82, -20, -128, 26, 82, 127, -106, -128, 66, 112, 65, -72, -2, 44, 17, -97, -128, 39, -24, 127, 3, -3, 41, -128, 109, 25, -27, 109, -5, -93, 34, -75, -6, 127, -128, -98, 9, 111, -20, 20, 125, 0, -128, 22, -13, -85, 37, 29, 26, -43, 119, -104, -31, 113, -55, 44, 83, -108, -128, 96, 49, -36, 10, -66, -66, 41, 114, -68, -44, 127, -2, 25, -12, 1, 112, -128, -41, 93, -128, 103, 76, -128, 87, 40, -128, 19, 76, -102, 74, 90, -128, 31, 100, -30, -41, -95, 121, 127, -128, -17, 117, -13, -116, 45, 115, 4, 19, -103, 3, -49, -64, 9, -48, 55, -38, 87, 87, -128, -15, 14, -86, 127, 23, -89, 30, 22, 25, -68, -20, 5, -36, 21, 127, -76, -47, 24, 27, 113, 11, -77, -97, -26, 125, 80, -42, -61, 18, 86, -61, -114, 36, 10, -26, -12, -88, 127, 27, -116, 70, 88, -99, 23, 19, -117, 48, 13, 20, -27, 70, 0, -97, 61, 25, -59, -11, 58, -9, -30, -38, 91, 123, -45, -128, 24, 82, -95, 52, 9, -119, 105, -43, -36, 127, 38, -107, -79, 45, 79, 52, -128, -108, 83, -37, 76, 127, -99, -64, 1, -19, 3, -34, 0, 3, 49, -29, 68, 72, -98, 109, -68, -128, 17, 112, -2, -115, 17, 11, 37, 124, -22, -106, -24, -30, 15, 93, 1, 6, -15, -20, -48, -8, 3, -69, 20, 104, 12, -35, -1, -58, 127, 119, -115, -82, -3, 7, 47, 38, 8, 24, -128, -10, 115, -100, 17, 104, -31, 17, 51, -94, 34, 91, -128, 47, 81, -128, 17, 62, -7, 58, 59, -128, 46, 90, 17, -66, -128, 111, 120, -113, -71, 127, 17, -19, -44, 14, -44, -20, 8, 14, 121, 9, 11, -127, -39, 127, -110, -128, 86, 122, -24, -128, 77, 110, -15, -49, 34, 59, -88, 61, -61, -12, 102, -90, 90, -94, -22, -8, -19, 70, 3, 83, -115, -34, -30, 92, 5, -128, 127, 58, -54, 44, -114, 37, 106, -127, 48, 66, -19, -108, -23, 127, -90, -30, -31, 21, 18, 6, -14, -22, 87, -128, 79, 48, -9, -46, -20, -1, -92, 19, 6, 63, 116, -102, -117, 127, 12, -49, 19, 14, 95, -128, 34, 81, -128, -11, 47, -30, -41, 55, -19, 29, 112, -78, -123, 127, 63, -28, -37, -95, -36, 42, 127, -2, -79, 12, -8, -34, -51, -56, 127, 18, -108, 38, 28, 106, -58, -28, -39, -76, 127, 72, -128, 58, -3, -81, 44, 10, 85, -17, 28, -14, -110, 74, 34, -128, -42, 126, 89, -100, -69, -25, -29, 1, 73, 12, -60, 54, -24, -13, 121, -46, -53, 127, -83, -97, 63, 91, -45, 12, 104, -128, -100, -1, 127, 127, -128, -81, 127, -4, -4, 11, -95, 81, -54, -128, 126, 17, -123, -11, 5, 127, 91, -82, -25, -85, 20, 97, -72, 51, 42, -102, 30, 80, 31, -28, -51, -24, 72, 34, -128, -107, 85, 82, 40, 69, -110, -57, 24, 14, -7, -59, 97, 92, -94, -128, -12, 127, -9, -127, 123, -38, -128, 127, 44, -82, 2, -10, 2, 13, 61, 12, -128, 1, 46, -105, 68, 57, 18, 51, -128, 69, 2, -18, 80, -124, -42, 25, 24, 74, 4, -62, 54, 0, -2, 69, -128, 17, 127, -128, -53, 18, 82, 43, -128, 73, -11, -55, 127, -128, -82, 44, 22, 90, 7, -28, -100, 11, 94, -29, 38, -37, -61, 96, -45, -54, 80, -109, 41, 127, -59, -120, 14, 127, -8, -51, -24, -43, 61, 46, -61, 69, 31, -29, -92, -93, 94, 54, 26, 3, -41, -85, -91, 3, 127, 105, -125, -57, 120, 117, -128, 2, -38, -78, 48, 27, -27, 58, -1, -85, 127, -86, 0, 6, -2, 112, -29, -128, 20, 127, -47, -35, 57, -54, -117, 60, 56, -123, 89, 99, -19, 2, -18, 45, -30, -20, -59, -48, 18, 98, -19, -123, 56, -4, -21, 10, 36, -52, -7, 124, 15, -128, 83, 42, -92, 41, 66, 0, -128, 127, 76, -62, 26, 47, -46, -117, -23, -48, 80, 23, 5, 115, -9, -40, -95, -78, 127, 115, -73, -128, 92, 25, -43, -8, 32, 9, -96, 123, 20, -29, -21, 37, -55, -120, 127, 13, -81, 107, 51, -128, 24, 120, -66, 71, -13, -35, -57, -13, -7, -40, 53, -27, 26, -62, 82, 127, -128, 4, 69, -115, -27, 80, 70, -107, -119, 107, 127, -63, -97, 87, 41, -91, 43, 119, -37, -128, -44, 127, -86, 1, 112, -51, -54, -22, 17, -18, 116, -47, -106, 126, -19, -90, 114, 73, -71, -40, -35, -89, 127, 117, -128, 90, -34, -96, 20, 11, -15, 27, 127, -128, -70, 4, 75, 102, -128, 68, -10, 27, -8, -105, 72, -91, 96, -34, -2, 15, -69, 22, -22, 106, -4, -69, -4, -59, 114, 39, -119, 120, 62, -128, -6, 53, 21, 7, -98, 127, 23, -128, 71, -1, 5, 83, -78, -1, 25, -9, 77, -49, -37, 1, -27, 105, -57, 17, 35, -51, -82, 71, 89, -128, 14, 32, -17, 4, -103, 127, 18, -124, -8, 98, 92, 3, -43, 14, -61, -71, 82, -61, -39, 62, 127, -3, -128, 15, 127, -11, -81, 30, 58, -126, 27, 48, 18, -53, -41, 5, -128, 114, 127, -4, -128, 15, 24, -39, 105, -105, 25, 68, -57, 4, 79, -54, -119, 79, 64, 3, -65, -57, 46, 25, -2, -9, -48, 23, 127, -58, -31, 116, -83, 5, -48, -108, 85, 44, 0, 6, 47, -29, 35, -12, -128, 55, 127, -44, -61, -57, 8, -21, 79, 0, -28, 127, -71, -114, -49, 35, 55, 45, 12, -110, 41, 120, -115, 65, 61, -128, 31, 64, -116, 127, 3, -128, 56, 79, 52, -88, 73, 15, -105, 92, 42, -121, 53, 115, -34, -31, -70, 91, -5, -111, 39, 122, -111, -109, 127, -43, -19, 70, 63, -96, 6, 29, -21, -37, 37, -31, 1, 21, -105, 79, -66, 82, -23, -97, 127, -11, 9, 19, -73, -26, 47, 26, -5, -56, 13, 75, -3, 43, -86, -92, -10, 19, 27, -1, 32, 20, -27, 24, -75, 25, 25, 13, 66, -21, -25, -97, 49, -12, -95, 127, 112, 24, -102, -79, 116, 31, -57, -40, -69, -25, -7, 127, 127, -75, -126, -79, 26, 10, 35, 14, 90, -7, 1, 42, -53, -111, 66, 87, -128, 93, 106, -89, -43, -46, 49, 127, -57, 37, 23, -128, 121, 21, -112, 3, -42, 65, -10, -3, 49, -10, -63, -40, 104, -62, 14, 106, -128, 35, 72, -9, 23, 36, 39, -49, -116, -98, 127, -29, -12, 53, -96, 73, -2, -73, 13, 87, -25, 5, 78, -53, -89, 32, 11, 6, 36, -21, 38, -87, -106, 87, 8, 86, 27, -31, -78, -23, 58, 15, 48, 7, -78, -2, 127, -11, -121, 59, 23, -128, 110, 73, -55, 43, -42, 3, -23, 74, -30, -14, 40, -83, 17, 70, 59, -37, -128, 48, 25, -43, 6, 9, 19, -81, 51, -42, 63, 127, -128, -8, 127, -2, -81, -96, 114, -75, -68, 127, -75, -88, 9, 92, 34, -65, -47, -85, 127, -3, -113, 31, -64, 105, 125, -104, 20, 15, -128, 53, 29, -42, 124, -25, -128, 8, -39, 127, -23, -26, 127, -102, -119, 57, 103, 22, -60, -66, 97, 78, -111, -106, 9, -63, 127, 89, -52, -115, 102, 1, -96, 102, 6, 30, -83, -35, 127, 0, -20, 6, -128, 71, 26, -96, 88, -69, 28, 126, -59, -32, 66, 42, -41, 21, -29, -128, 38, 79, -105, 65, 116, -56, 11, -94, -105, 73, 57, 37, 41, -19, -128, 31, 127, -113, -30, 70, -128, -2, 127, 25, -95, 58, -18, -105, 56, 110, -52, 19, -52, -42, 127, -128, -62, 97, -28, 79, -19, -108, 41, -60, 0, 9, 114, 70, 13, -95, -128, 108, 103, -116, 14, 82, -48, -7, -38, -21, 30, 116, 8, -25, -5, 37, -117, -96, 20, 7, 126, 69, 13, -128, -4, 57, -45, -7, 49, 32, 14, 72, -89, -61, -3, 94, -17, -128, 22, 127, -70, -63, 8, 11, 70, -105, 61, 127, -86, -54, -54, 75, 31, 2, -31, -10, 96, -58, -93, -46, 127, -3, -128, 47, 127, -42, -59, 71, -13, 45, -65, -19, 115, -128, 7, 127, -128, -5, 15, -76, 104, 41, -21, -39, -32, -21, 59, -34, -98, 14, 94, 56, 24, -66, -107, 127, -104, 8, 92, -128, 127, 110, -66, -92, -104, 127, 106, -28, -7, -128, 59, 0, 14, -22, -19, 127, -46, 0, -59, -25, 0, 11, 54, -17, -35, 4, 8, 66, -56, 0, 32, -22, 23, -1, -65, 40, 117, -73, -69, -39, 114, -64, -13, 36, -128, 103, 0, -52, -27, 68, 70, -112, 92, 57, -72, 11, -71, -93, 127, 58, -128, 127, 13, -128, 127, 77, -128, -21, 68, -46, -28, 42, 61, 105, 37, -99, -17, -41, -81, 0, 65, 89, -108, 48, 127, -22, -30, 9, -128, 18, 127, -128, -114, 117, 44, -81, 45, -31, -57, 27, 74, -15, -112, -4, 99, -8, -28, 12, -106, 60, 127, 7, -92, -28, 17, -9, 6, 111, -51, -19, 0, -74, 15, 109, -46, -100, 114, 37, -94, -47, 83, -59, -73, 34, 77, 71, 10, -128, 39, 127, -128, -112, 98, -32, 46, 83, -36, -47, -1, 115, -35, -30, 0, -103, 17, 127, -56, 29, -35, -128, 103, -49, -78, 49, 123, -58, -98, 127, -72, -120, 107, 103, -53, -44, -79, 5, 127, 3, -40, 17, -58, -128, 73, 57, -65, -12, 14, -9, 78, 89, -128, 74, 15, -52, 2, -37, 127, -112, -96, 31, 23, 120, 100, -63, 13, -88, 8, 49, -8, -85, -3, 45, -110, 37, 107, 5, -106, -15, -30, 6, 71, 90, -6, -56, 18, -40, -80, 65, 88, 74, -103, -128, 60, -61, 124, 47, -128, -12, 88, 34, 15, 49, -96, -113, 115, 127, -128, -49, 15, 70, -20, 26, 127, -128, 24, 44, -65, 74, -37, -15, 83, -100, 15, 127, -123, -22, 68, -30, -7, -77, -95, 127, 124, -23, -62, 4, -22, 1, 47, 9, -25, -45, -28, -26, 17, 41, -69, 32, 127, -128, -98, 88, 6, -23, 78, -60, -80, 8, 90, -15, -55, 47, -71, 0, 9, 68, 61, -94, 32, 127, -128, -128, 127, 9, -49, 99, -113, -43, 64, -39, 76, 53, -128, 58, 127, -80, -42, -91, 91, 31, -77, 2, -64, 115, -24, -18, 72, 0, -87, 30, 74, -128, -23, 127, 29, -83, -13, 7, 34, 1, 2, 4, -48, -64, 127, -27, -22, 125, -128, 29, -2, -128, 100, 104, -30, -92, -26, -14, 100, 55, -62, -12, 39, -51, -48, 111, -60, -29, 114, -37, 48, 0, -128, 97, 103, -48, 48, -14, -43, 44, -73, 13, -17, -97, -19, 127, -7, -128, 24, 21, -18, 40, 127, -65, -104, 6, -59, 127, 40, -128, 103, 70, -40, 82, -76, -126, 34, 94, 29, -17, 47, -47, -128, 127, -7, -98, 64, -22, -15, 30, 15, -13, -56, 39, 127, -15, -98, -8, 40, 44, -66, -77, 78, 48, 78, -66, -97, 46, -18, -70, -18, 58, 127, -74, -15, 48, -40, 8, 7, -27, -89, 86, -47, 73, -37, -26, 127, -112, 56, 11, -128, 55, -19, 58, 92, -128, 76, 127, -112, -128, 42, 106, -24, -76, 17, 92, 83, -120, -60, 19, -70, 24, -10, 68, 82, -128, 71, 61, -83, 74, 22, -81, 42, -4, -73, 127, -5, -128, -29, 110, 87, -105, 6, 45, -128, 88, 92, -128, 57, 24, -88, 127, 44, -60, 76, -103, -39, 108, 5, 74, -128, -28, 66, -41, 107, -42, -97, -11, -58, 110, 127, -128, -62, 127, -106, -75, 127, 65, -122, -72, 31, -27, -22, 57, 127, -106, -128, 83, 127, 7, -25, 58, -106, -128, 48, 105, 12, -108, 75, 86, 9, -68, -72, 116, -87, -62, 91, -64, -62, 121, 37, -120, 17, 44, -12, 105, 0, -128, 59, -5, -23, 127, -75, 14, 46, -85, -72, 90, 37, -96, -6, -74, 116, -23, -1, 127, -108, 30, 52, -70, -112, -1, 65, 30, 125, -128, -15, 111, -105, 90, -74, -37, -10, 14, 117, -68, -86, 46, 119, 43, -128, -49, 127, -35, -91, -62, 81, 43, 57, -73, -71, 61, 2, -35, -13, 58, -108, 87, 127, -128, 22, 81, 12, -62, -38, 120, -61, 22, -65, -119, -2, 61, 122, -4, -17, -23, -68, 77, -38, -110, 23, -25, 102, 43, -47, -15, 15, 36, -87, -2, 78, -76, 81, 127, -128, -97, 127, 75, -91, -93, -12, 127, -108, -15, 127, -128, -64, 45, -59, 63, 62, 3, 6, -60, 12, -45, 62, 112, -62, 32, -99, 18, -7, -63, 96, -79, 108, -4, 12, 4, -73, 127, -128, 59, 39, -128, 127, 56, -128, 70, 21, -128, 25, 61, 61, 14, 86, -128, -25, 111, 8, -18, 4, 27, -38, -27, 32, 28, -66, -36, 51, 59, -24, -62, -30, -1, 3, 11, -10, 86, -74, -12, 110, -35, 12, -44, -71, -25, -11, -12, 73, 97, -7, -73, 35, 127, -128, 6, 97, -34, 72, -79, -18, -83, 61, 72, -13, -36, -104, 0, 68, 122, -128, 26, 126, -27, 15, -128, 23, 12, -87, 55, -40, -1, 92, 93, -107, -128, 107, 12, -38, 125, 11, -123, 55, 41, -128, 28, 55, -66, 81, -47, -31, 113, 22, -46, 62, -39, -25, 0, 28, 20, -128, 122, 40, -96, -78, 86, 44, 35, -15, -128, 121, 127, -114, 0, 54, -116, -73, 120, 0, 71, -38, -38, 127, -128, -78, 56, 68, -47, -42, -30, 108, 2, -93, 86, -81, -22, 122, -28, 22, 8, -128, 113, 26, -128, -5, 127, -12, -92, 97, -36, -2, -18, -106, 127, -23, -128, 20, 7, 127, -20, -13, 49, -46, 72, -87, -4, 121, -127, -13, 127, -75, -82, -15, 77, -25, -49, 114, -68, -120, 56, 58, -7, -40, 58, 39, 23, -42, -119, -10, 98, 99, -57, 3, 63, -90, -64, 28, -48, 65, 25, -76, 59, 88, -49, -47, -45, 93, 107, -60, -49, -73, 124, -40, -65, 58, 42, 3, -128, 53, -35, -81, 116, 24, -5, 68, -94, -86, 127, 45, -68, 32, 82, -107, -21, 87, -128, 76, 127, -128, 30, 68, 15, -51, -92, 103, 61, 24, -80, -66, -75, 88, 47, -128, -3, -8, 39, 112, 13, -119, -44, 127, 23, -79, 29, -5, -108, 62, 127, -52, -95, -55, -27, 99, 88, -10, -119, -19, 127, 53, -46, -60, -29, -47, -1, -14, -31, 66, 0, -49, 99, -75, 63, 127, -128, -21, -51, -46, 112, 54, -17, 12, -56, 5, 81, -128, 66, 127, -119, 63, -44, -128, 127, -35, -56, 5, -41, 127, -15, -46, -53, -68, 54, 34, 73, 12, -77, -57, 53, 86, 24, 13, -86, 7, 65, -20, -90, -15, 127, -76, -81, -57, 103, 28, -102, 120, 31, -21, -127, 43, 96, -30, -3, 24, 0, -92, -88, 102, 102, -95, -23, -71, 95, -15, -14, 110, -100, -51, -51, 83, 36, 45, -42, 25, 21, -42, -35, -8, 127, -70, -80, 53, -47, -37, 31, 51, 95, -92, -98, 122, -23, -107, 0, 44, 72, -2, 0, 65, -52, -58, 29, -60, -31, 85, -70, -78, 127, -76, 7, 0, 15, -8, -21, 127, -128, -81, 127, -82, -70, 127, -29, 41, -48, -82, -4, 58, 65, -25, 38, -47, -19, 28, -93, -5, 110, -68, -112, 108, 53, 15, 58, -128, -8, 81, -74, -42, 89, -29, -54, 27, -18, 107, -87, 15, 127, -95, 27, 91, -128, -92, 86, 71, 53, -122, -71, 122, -10, -22, 72, -61, -29, 22, -49, -12, 114, 18, -48, -31, 29, 24, -2, 87, -36, 4, -25, -128, -40, -9, 124, 76, -128, 94, -9, 6, 0, -63, 58, 28, -12, -76, 127, 57, 8, -73, -73, 91, -8, 5, 0, -103, -31, 107, 98, -77, -3, 36, -128, -61, -4, 127, 111, -128, -66, 127, 53, -108, -108, 39, 28, -12, -44, 114, 10, -128, 87, -58, 78, 127, -86, -112, -31, -30, 127, -8, -82, 127, -106, -128, 127, 7, -76, 115, 39, -128, -4, 127, -128, -128, 90, 77, -44, 91, -29, 5, 9, -128, 79, 29, -85, 110, 52, -38, 6, 52, 62, -6, -29, -92, -3, -37, 59, 127, -30, -128, -4, 114, -21, -92, -96, 106, 87, -39, -6, -59, 63, 47, -81, 62, -56, -41, 127, 2, -102, 5, 3, 58, 57, -128, 34, 54, -128, 95, 89, -128, 22, 60, 18, 87, -128, 30, 105, -25, -94, 25, -17, -87, 127, 59, -93, -106, 127, -65, -114, 51, 27, 9, -68, 10, 97, 44, -105, -66, 127, -28, -70, 34, 47, 74, -21, -62, -48, 94, 61, -71, -78, 76, -20, -12, 48, 44, -128, -54, 127, -87, -128, 56, 93, 30, -57, 25, 77, -106, -9, 102, -109, 12, 29, -128, 123, 127, -128, -87, 69, 3, 79, 1, -98, 14, -27, -2, -8, 40, 127, -21, -128, -40, -11, 112, 9, -37, 127, -76, -109, 0, 55, 102, -122, -71, 127, -102, 43, 127, -128, -3, 127, -79, -15, -48, -93, 44, 61, 90, -2, -49, 85, -107, -114, 73, 73, 71, -120, -128, 69, 124, -31, -47, 95, 89, -128, -95, 28, -46, 127, -27, -83, 108, 48, -125, 58, 97, -128, -4, 10, -68, 5, 127, -6, -45, 20, -10, 51, -31, 52, 69, -76, -119, 52, 127, -36, -77, -53, -86, 127, 72, -56, 80, -103, -128, 25, -27, 123, 127, -29, -87, -17, -45, -17, 127, -44, -99, 64, -12, 76, -31, -31, 11, -124, -8, -26, 122, 127, -7, -128, 28, 127, -60, -37, -10, 4, 0, -10, -36, 0, -81, 108, 83, -74, 6, -38, 5, 0, 78, -78, -19, 116, -127, 32, 93, -105, -58, 89, 75, 51, -74, -86, 13, -15, -23, -56, 21, 78, 83, -32, -121, 28, 19, -14, 82, 61, 28, -120, -128, 39, 3, -24, 90, 119, -107, 37, 26, 3, -81, -61, 127, -128, 23, 122, -128, 72, 28, -1, 39, -68, 78, 39, 10, -97, 12, 81, -95, -3, -4, 2, 6, -93, 49, 111, -17, -98, 11, 108, -12, -122, 22, 80, -128, 85, 31, -128, -1, 127, -22, -128, 124, 47, -65, 85, 58, -20, 29, -128, -8, 127, -27, -111, 57, 107, 4, -59, -71, 93, 5, -51, -37, -11, 9, 38, -6, 4, 85, -3, -83, 6, -10, -45, 41, -21, 52, 52, -108, 54, -6, -43, 39, -58, -61, 126, -3, -128, 91, 59, -90, 82, 83, -128, 108, -15, -102, 127, -121, -56, 96, -128, 66, 125, -128, 32, 6, 59, -24, -128, 127, -35, -1, 71, -63, -79, -47, 127, -81, -117, 127, -65, -75, 1, -60, 10, 35, 89, 4, -96, 97, -11, -128, 127, -61, -13, 127, -128, -23, 127, -128, -11, 120, -76, -102, 126, -34, -61, 127, -5, -107, -56, 127, 51, -57, 48, -55, -69, 9, 104, -82, -128, 119, 103, 49, -119, -99, 44, -19, -3, 90, -34, 32, 87, -29, 15, -70, 66, -11, -128, 99, 46, -8, 99, -128, -19, 24, -128, 116, -7, -55, 94, -23, -80, 122, 7, -116, 25, 21, 102, -47, -36, 5, -12, -44, 11, -14, -3, 127, 0, -95, -44, 26, 85, 71, -40, -82, -100, -27, 110, 114, -32, -128, 34, 94, -110, 62, -35, 54, 9, -59, 14, -59, 17, -61, 48, 62, 79, 53, -128, -80, 117, 91, -102, -112, 90, -9, -46, -11, 105, -46, 19, 114, -52, -32, -74, 40, 6, 77, -24, -7, 56, -21, -58, -9, 27, -93, -55, 127, -46, -15, 57, -55, -17, 36, 124, -128, 45, 56, -85, 127, -36, -75, 77, -27, -63, -5, -46, -36, -10, 69, 53, -91, 45, 127, -79, -104, -9, 81, 71, 10, 9, -126, 43, 127, -125, -62, 13, -91, 127, 110, -96, -18, 58, 30, -128, -37, 66, 25, 53, -86, 19, -4, 40, -30, -56, 127, -95, 41, -27, -65, 37, 21, 68, -66, -49, -53, 0, 55, 55, -9, -78, 29, 65, 51, -15, -12, -70, -44, 68, 43, -22, -109, 85, -45, -41, 41, -88, 85, 36, -105, 115, 66, -128, -68, 121, 127, -128, -71, 34, -59, 72, 26, 32, -45, 0, 20, 7, 24, -57, 127, -100, -57, 117, -104, 11, 127, -55, -59, -3, 90, -17, -21, 25, -108, 78, 10, 22, 32, -100, -9, 45, -63, 75, 4, -58, 116, -114, -113, 78, -18, 87, -19, -40, 42, 40, 28, -45, -21, -122, 71, 81, -35, -14, 30, -92, 43, 41, -128, 127, 95, -38, 23, -107, -69, 56, 110, 68, -128, -105, 109, -43, -99, 127, 78, -79, -70, 2, -21, -11, 127, -79, -128, 127, 78, 23, -128, 24, 64, -82, -27, 78, 25, -107, 32, -27, 110, -63, -31, 127, -104, -66, -10, 21, 115, -78, -44, 75, -35, -53, 0, 10, 112, 9, 7, -54, -126, 110, -8, -8, -38, -9, 46, -46, 57, 80, 22, -91, 17, 24, -69, -11, -11, -2, 9, -41, 82, 21, -68, -64, 114, 39, -46, 62, -76, 46, 55, 36, -128, -112, 42, 23, -14, 122, -4, -128, 1, 113, 10, -128, 127, 9, -44, 127, -45, -89, -110, 55, 0, 97, 24, -20, 1, -128, 98, -35, 35, 55, -100, 30, 122, -59, 0, 34, -52, 65, 7, 15, -66, -65, 37, 106, -75, -49, 119, -58, -107, 127, 8, -93, 82, 5, -51, -31, -7, 114, -47, -77, 97, -102, -54, 127, -49, -93, 12, 3, 85, -70, 39, -5, -13, 8, -116, 127, 30, -126, 124, -30, -119, 93, -25, -66, 32, 42, 54, -22, 0, 121, -125, -99, 127, 42, -23, 7, -88, -95, 79, 74, 44, -71, 6, 12, -128, -31, 100, 127, -66, -98, 28, -45, 72, 100, -123, 12, -27, 64, 51, -28, 41, -34, -109, -82, 127, 127, -121, 36, -52, -78, 127, -76, -94, -34, 96, 3, -104, 3, 103, 54, -10, 57, -89, 29, -51, -115, 127, -47, -60, 127, 7, -73, -63, -11, 79, -52, -12, 63, -128, 112, 70, -6, -91, 6, 98, -122, 12, -20, -56, -21, 127, 45, -119, -9, 87, 72, -49, 77, -94, -128, 127, 65, -81, 24, -116, -1, 122, -69, -89, 95, 18, -20, 3, -28, -35, 26, 127, -128, -1, 127, -128, 14, 36, 19, -4, -39, 127, -128, -64, 127, -2, -75, 12, -47, 58, 127, -128, -115, 49, 71, 80, -90, -75, 32, 41, 36, 1, -53, -72, -6, 125, 121, -17, -77, -117, 54, 52, -71, 24, 34, 74, -85, 37, 6, -110, 83, -49, 23, 9, 46, 48, -103, -5, 53, 60, -28, -32, 92, -99, 30, 19, -128, 93, 14, -123, 49, 25, -99, 117, 127, -77, -128, 23, 127, -79, -128, 116, 115, -26, -107, 45, 92, -53, 37, -128, -5, 127, -54, 42, 42, 12, -87, -102, 25, 21, 83, -28, -60, 35, 49, 28, -4, 41, -116, -128, 127, 15, -19, 41, -113, 25, 51, -34, 63, -102, 20, 127, -47, -44, 7, -44, 27, -42, -3, 63, -128, 25, 43, -34, 115, 9, -70, 69, 42, -110, -5, -40, -1, 45, -55, 107, 43, -46, -5, -91, 25, 127, -48, -72, 94, -1, -64, -81, -30, 4, 4, 85, 2, 11, 7, -96, 47, 10, -8, -4, -100, 1, 100, -34, 34, -1, 17, 61, -128, 25, 59, 100, 10, -128, 26, 95, 6, -39, -105, 11, 127, 28, -106, -77, -1, 65, -26, -37, 77, -27, 25, -58, 70, 31, -29, 95, -128, 22, 64, -128, 82, 127, -66, 21, -64, -39, 70, -53, 19, -22, -106, 2, 127, 40, -23, 45, 0, -27, -99, -44, 103, 48, -52, -126, 70, 96, 0, 2, -77, -3, -24, 0, 88, 5, -94, 69, -75, -32, 127, -81, -111, 7, 68, 61, 39, -116, 4, 127, -42, -30, 11, -102, 2, 26, -39, -9, 36, 18, 11, 39, -128, 22, 0, -13, -10, 7, 124, -8, -107, -6, 119, 53, -110, -114, 6, 108, 0, -26, -5, -62, 75, 127, -62, -47, -57, -37, 111, -81, -46, 48, 47, -1, -66, 65, 40, -69, 38, -29, -80, 11, 127, -57, -17, 127, -128, -128, 59, 91, -26, 66, -25, -128, 127, 92, -27, -59, -9, 4, 35, -14, -86, 56, -35, 2, 105, -7, -71, 64, 58, -11, -54, -80, -65, -28, 127, 27, -104, 56, 127, -128, -17, 51, -128, 36, 58, 85, 35, 32, -127, 28, -22, -87, 85, 45, -55, -128, 126, 20, -110, 11, 127, -43, 6, 46, -128, 127, 127, -53, -114, 36, 51, -62, -57, 63, 112, -128, -13, 81, -66, -34, 79, -57, -85, 127, 57, -94, -17, -37, 120, -37, -41, 127, -128, -45, -14, 8, 127, -114, -13, 103, -27, 5, -81, 6, 47, -103, -58, 5, 41, -12, 108, 18, -20, 44, -28, 41, -123, -88, 8, -5, 127, 79, 9, -87, -18, 23, -87, 35, 60, -77, 17, -18, -41, 21, -64, 93, -27, -41, -30, 127, 121, -29, 3, -121, 21, 99, -25, -85, -96, 105, 70, -80, -10, 4, -61, 100, 120, -73, 7, -75, -1, 127, -61, -128, 79, 26, -79, 52, 0, 7, -10, 5, 61, -102, -86, 127, 100, -11, -128, 47, 56, -23, 91, -19, 5, 22, 15, -128, 53, 58, -89, -38, 26, 25, -109, 127, 85, -116, 17, 107, 6, -59, 2, 3, -61, 66, 21, -91, -65, 53, 24, 65, -69, -69, 72, 9, 92, 18, -128, 14, 96, 7, -76, -105, 11, 112, 51, -128, 98, 1, -96, 44, -44, 72, 39, 24, 72, -46, 0, -11, -108, 9, 104, -83, -26, -6, 11, 64, -10, -23, -95, 53, 38, 49, 8, -25, 9, -10, -19, -55, 37, 3, 70, 30, -128, 4, 127, 6, -128, -62, 108, -54, -37, 27, -44, 37, 127, -49, -27, 41, -128, -5, -1, 39, -26, 93, 71, -128, 119, -14, 14, 77, -128, 23, 32, -46, 119, 13, -24, 11, -22, -47, -90, 49, 29, -43, -30, 41, -29, 19, 4, -56, 116, 36, -102, 81, -11, 57, 19, -128, 17, 1, 80, 39, 35, -59, -128, 53, 127, -76, -128, 127, 121, -128, -80, 113, 45, -103, -85, 127, 127, -5, -19, -51, -13, -34, -64, 111, -39, -115, 17, 6, 71, 32, 35, -66, -93, 53, -1, -24, 48, 96, -23, -109, -27, 127, 14, -40, -74, 15, 44, 41, -47, -46, 77, -22, 53, -75, -42, 97, 96, -128, 4, 127, -128, 23, 90, 3, -36, -74, 79, -102, -60, 124, -48, 45, 27, -102, 77, 81, 6, -128, 31, 56, -60, -56, 30, -19, 74, 20, -35, 74, -87, 76, -72, -114, 127, 116, -120, -77, -21, 81, 127, -128, -70, 63, -30, 46, 98, -44, -96, 45, -63, -78, -1, 93, 125, 30, -128, -125, 127, -38, -31, 81, 31, 71, -56, -3, 28, -89, 35, -42, -39, 111, -54, 11, 113, -28, -81, 34, 62, -128, 29, 127, -111, -108, 64, 82, -119, 25, 85, -109, 48, 92, -55, 51, -21, -19, 14, -128, 121, -31, 14, 6, -25, 12, -20, 14, -128, 124, 122, 45, -128, 19, 26, -128, -3, 35, 6, 74, 127, -1, -64, -91, 10, 69, -65, 47, -25, -52, -26, 70, -14, -23, 127, -34, -61, -102, -22, 107, -37, -123, 127, -37, -25, 78, -104, -22, 7, 40, 0, 13, 1, 24, -17, 62, 3, -128, 127, -35, -61, 43, -15, 45, -12, -25, -28, 78, -54, -102, 127, 114, -128, -25, 127, -68, -45, -19, -56, 113, 1, -2, -32, -35, 39, -21, 77, -37, -28, 40, 69, -81, -44, 73, -82, 57, -36, -117, 63, 41, 59, 70, 7, -62, -128, 87, 94, -128, 110, 26, -73, 94, 39, -128, -10, 19, -14, 110, 43, -88, -128, 36, 53, -39, 77, 23, -47, -7, -8, 96, 11, -59, 39, -97, 42, 113, -18, -46, -27, -13, -31, 80, 51, 2, -128, 100, 45, -75, 58, -128, 97, 78, -64, -52, -58, 127, 11, 32, -77, -98, 49, 43, -37, -105, 41, -2, 6, 127, 32, -69, -17, -77, 44, 127, -13, -73, 3, -81, -60, 127, 103, -128, -66, 127, -119, -90, 107, 85, -2, -57, -59, -77, 127, 11, -126, 1, 29, 28, 19, 71, -47, -117, 106, 113, -14, 12, -115, -58, -13, 90, 73, -28, 70, -128, -69, -13, 17, 110, 40, 17, 11, -113, -28, 86, -62, -53, 75, 104, -15, -115, 59, 32, -88, -53, 57, -32, -20, 28, -3, 120, -22, 34, -31, -128, 115, 127, -99, -26, -71, 51, 8, 24, 72, -63, -39, 56, -63, -53, 82, -93, -8, 23, 17, -10, 13, -4, -26, 39, 17, -32, -24, 20, 15, 102, -39, -107, 122, -19, -95, 23, -12, -26, 47, 127, -37, -127, -20, 48, 58, 66, -15, -107, -9, 23, 44, 61, 31, -114, -51, 44, -28, 43, 43, -93, 6, -8, -14, 68, 12, 46, 48, -14, -57, -92, -7, 96, 99, -128, -128, 65, 94, 69, 12, -122, -69, 63, -37, -6, 12, -2, -71, 127, 15, -128, 127, 2, -128, 92, -44, 75, 82, -37, -36, -17, 75, -45, 20, -43, 12, -55, 71, 0, -60, 127, -128, -26, -3, 74, 64, -85, 31, -30, 4, 40, -4, 49, -103, -11, 21, 22, 127, -10, -93, -128, 105, -11, -87, 127, 64, -48, -112, -64, 13, 32, 89, 37, -114, 24, 106, -72, -44, 31, 52, 43, 44, -110, 17, 14, -123, -47, 106, 10, -104, 52, 78, 15, -100, 49, 35, 12, 40, -82, 39, -63, -122, 92, 3, 46, 13, -128, 120, 127, -128, -120, 111, 124, -128, -128, 3, 117, 40, -10, 70, -8, 3, -88, -1, -5, -98, 44, -27, 11, 127, -15, -128, -18, 127, -20, -128, 43, 115, 79, -85, -52, 102, 0, -57, -12, 22, 63, -59, -28, 90, -128, -36, 127, -76, 55, 61, -27, 66, -5, -128, -18, 120, 14, -23, 6, -76, -46, 0, 12, 105, 26, -71, 47, -54, -79, 22, -13, 42, -32, -9, 19, -48, 12, 30, 109, -24, -58, 25, -109, 80, 47, 18, 70, -128, -44, 127, -75, -45, 57, 37, -47, 24, -39, -6, 38, 26, 28, -128, 27, -31, 65, 127, -128, 5, 24, -66, 74, 42, -40, -98, 74, 81, -46, -58, 120, -63, -93, 127, -14, -30, 34, 73, -89, -115, 32, -52, 41, 127, 25, -26, -13, 40, -105, 4, 102, -106, -1, -14, -6, 42, -60, 77, 126, -15, -128, -26, 86, -17, -97, 12, 31, 57, 66, -79, 32, -77, -80, 31, 114, 88, -128, 56, 2, -59, 97, -1, -96, 52, 127, -128, -23, 127, -128, -48, 127, -4, -128, 2, 127, -102, -113, 127, 15, -128, 51, 105, -80, 13, 34, -128, 26, 111, -26, -15, -21, -47, 56, -10, 42, 23, -23, -11, -83, 102, 45, -52, 85, -80, -52, 76, -114, -5, 127, -56, -128, 82, -21, -98, 18, 127, -1, -23, -21, -64, 127, -42, -110, 0, 53, -35, 72, 1, -126, 127, 13, -112, 29, -27, -57, 127, 31, -128, 127, 65, -111, 38, -26, -95, 127, -29, -63, 27, -110, 24, 127, 78, -37, -32, 5, 35, -69, -106, 127, 64, -110, -7, 80, -29, -31, 80, -73, -57, 127, -9, -128, 99, 73, -51, -39, 11, -25, -46, 83, 127, -114, -65, 70, -27, 23, -80, 108, 127, -108, -35, 37, -66, 66, 12, -128, -56, 95, 100, -92, -83, 98, 103, -54, -36, -26, 72, -49, -128, 127, 93, -128, 51, 62, -61, -86, 69, 9, -8, 71, -128, -4, 44, 90, -56, 41, 54, -128, 123, 127, -114, -105, 121, -69, -26, 40, -128, 127, 78, -128, 73, 127, -88, -29, -75, 64, 104, -128, -35, -52, 127, 29, -82, 46, 54, 40, -128, -92, 127, -39, -46, 115, -68, -22, -57, 43, 68, 26, -97, 15, 10, 26, 48, -63, 80, 39, -31, -123, -82, 127, 66, -128, -8, 105, 24, 64, -93, -109, 104, -41, -88, 127, 25, -128, 120, 122, -115, 51, -54, -72, 11, 82, 108, -117, -60, 2, 86, 117, -128, -27, 27, 32, 46, -98, 92, 43, -128, 43, 37, 0, -14, -79, 44, 38, -68, 1, 122, -85, 17, 27, -68, -47, -63, 59, -30, 47, 104, -115, -6, 96, 22, -73, -20, 93, 31, 20, -105, -128, 127, -12, -62, 70, 47, -14, -102, 44, 61, -9, 0, 6, -61, -3, -41, 22, 122, -128, -42, 99, 52, -52, 6, 0, -80, -7, 47, 114, -93, -48, 117, 68, -128, -1, 27, 15, 49, -10, -20, 2, -55, -24, 97, -64, 39, -6, -128, 68, 127, 7, -102, 2, 14, -12, 6, -47, 11, -95, 105, -24, 28, 2, -104, 127, 72, -55, -55, -82, 17, 28, -69, 17, 7, -21, 114, 37, -128, 95, 26, -32, 122, -60, -97, 93, -48, 2, 125, -19, -102, -19, 27, -46, 79, 43, 20, -65, -4, 14, -86, 12, -72, 96, 73, -91, -76, 68, 98, -128, -5, 127, 49, -128, 10, -19, 48, 79, -128, -35, 102, 127, -81, 6, 72, -127, -61, 127, -58, 6, 4, -96, 127, -102, -113, 106, 107, -88, -38, 93, -34, 2, 49, -87, -114, 40, 116, 98, -119, -92, -1, -29, 122, -4, -22, 8, 24, 69, -55, 43, -13, -54, -9, -21, -36, 66, -37, -5, 127, -60, -17, 111, -123, -32, 61, 5, -37, -34, -17, -7, 127, -17, -8, -103, -37, 127, -22, 28, 0, -61, -21, -34, 32, 15, 14, -59, 1, 93, 12, -15, -40, -90, -41, 8, 75, 127, -64, 5, 92, -128, 34, 112, -128, -107, 127, 99, -26, -128, -22, 85, 10, -85, 8, 28, -12, 127, 18, -62, -107, -70, 80, -7, 56, 95, -20, -15, -76, 34, -38, -79, 39, 4, 109, -25, -51, 20, 43, -58, -96, 85, -41, -77, 100, 91, -49, -83, -23, 127, -91, -61, 127, 42, -117, 0, -24, -112, 71, 90, -61, -124, 117, 72, -106, -29, 35, 53, -10, -71, 56, -40, 36, 127, -7, -128, 28, -31, 10, 126, -76, -105, 48, 109, -90, 6, -59, 43, 20, -128, 127, -36, -57, 127, -7, -125, -94, 108, 43, -128, 32, 81, -23, -5, -17, 74, 71, -128, 29, 81, -128, 120, 59, -119, -60, 66, 49, -44, 49, 82, -70, -128, 92, 113, -21, -57, -82, 39, 58, -11, -26, 61, -12, -128, 95, 127, 23, -99, -77, 30, -55, 15, -45, 86, 113, -128, 94, -56, -62, 90, -14, 68, -111, 10, 28, -114, 127, 45, -32, 27, -49, -90, 65, 99, -4, -21, 1, -20, -127, -59, 102, -27, 35, 122, -128, 92, 18, 11, -21, -128, 85, 46, -19, -30, 57, -96, 46, 122, -128, 73, 17, -128, 23, 127, -80, 38, 52, -128, 127, 26, -12, -37, -83, 104, 43, -68, -98, -7, 127, -49, -103, 110, 41, 17, -31, 12, -93, -98, 127, 36, -97, 36, 69, -110, 28, 80, -46, 66, -92, -69, 95, -32, 48, 108, -34, -8, -106, -44, 94, -103, 20, -3, 2, 127, -70, -69, -6, -80, 37, 10, 63, 93, -22, -82, -78, 127, 43, -124, 2, -60, 53, 71, -87, -81, 127, 127, -128, -47, 119, -25, 9, 41, -11, -60, -32, 57, -73, -13, 95, 2, -97, 42, 18, -112, 111, 76, -13, 59, -128, -10, 117, -96, -25, -65, 80, -4, -40, 83, -92, 107, 35, -128, 49, 123, -51, -63, 64, -36, 32, 114, -2, -65, -42, 19, 65, -63, -52, 55, -45, -66, 94, 18, -128, 95, 127, -76, -95, 61, -69, 4, 127, -19, -128, -58, 127, 102, -71, -15, -18, -128, 63, 127, -115, -103, 62, 90, -26, 7, 34, -128, 22, -23, -21, 117, -28, -128, 107, 24, -74, 108, -22, 39, -43, -90, 88, 78, -72, 14, 38, -114, 15, 127, -71, -119, 7, 32, 1, 15, 127, -30, -56, -25, -91, 39, 121, 21, -107, -1, -2, -13, -5, 61, 22, -102, 108, 34, 12, -44, -46, -35, -93, 95, 75, -5, -63, -91, 127, 2, -36, 34, 28, -8, -107, -23, -43, 127, 21, -60, -5, -61, -34, 55, 127, -53, -105, 108, -107, 20, 127, -128, 65, 43, -28, -41, 0, 7, 42, -40, 1, 92, -12, -91, -76, 23, 102, 19, -120, 10, 61, 90, -99, -7, 92, -45, -82, -38, 127, -35, 3, 66, -53, -65, -113, 127, 87, -128, 83, 17, -61, 80, -26, 7, 64, -53, -95, 85, -11, -95, 96, -47, 2, 127, -119, -120, 77, 31, 51, 85, -98, -76, 80, 38, -65, 42, 54, -71, -25, 57, 30, -128, -103, 18, 127, -52, -68, 127, 0, -103, 3, -60, 48, 99, -128, 120, 71, -62, 81, -97, -91, 107, -23, -71, 8, 39, 53, -75, 88, -49, 5, 80, -85, 4, -98, 88, 94, -88, -13, -38, 58, 56, 6, -52, 0, 77, -86, 74, -52, -109, 127, -2, -128, 65, 39, 4, -11, -30, 30, -96, -41, 75, -37, 51, 27, -22, 37, 0, 27, -53, 75, -59, -128, 27, 54, 13, 9, 64, 62, -128, -97, 122, -38, -22, 127, -103, -74, 127, -39, -35, -4, 36, 7, -95, 4, 111, -47, -73, 54, 32, -43, -79, 1, 120, 46, -128, 31, 3, -37, 98, -60, 9, -2, -98, 127, 47, -128, -5, 80, -51, 14, 38, -69, 71, -38, -30, 100, 26, -87, -91, 94, 47, 89, -97, -85, 113, 35, -22, -124, 29, -9, -13, 127, -91, -37, 60, 9, -47, 17, 124, -15, -128, -72, 20, 39, 58, -14, -54, -35, 61, 49, -98, 76, 103, -29, -69, -70, -34, 121, 15, -128, -3, 64, 127, -7, -102, -42, -51, -31, 127, -57, -8, 27, -6, 108, -44, -27, -4, -34, -90, 69, 72, -117, 8, 127, 30, -39, -3, -45, 43, 29, -44, -95, -21, 19, 22, 126, -5, -128, 14, 103, 23, -74, -91, -39, 121, -15, -80, 127, 35, -60, -73, -70, 87, 54);
    constant SCENARIO_ADDRESS2 : integer := 25000;    -- This value may arbitrarily change
  
    constant SCENARIO_LENGTH3 : integer := 47;
    constant SCENARIO_LENGTH_STL3 : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH3, 16));
    type scenario_type3 is array (0 to SCENARIO_LENGTH3-1) of integer;
    signal scenario_config3 : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL3(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL3(7 downto 0))),    -- K2
                                                      127,                                                        -- S
                                                      -1, -1, 8, 0, -8, 1, 1, 1, -9, 45, 0, -45, 9, -1           -- C1-C14
                                                      );
    signal scenario_input3 : scenario_type3 := (-115, 60, -102, 14, -112, 7, -68, -122, -96, 120, 8, -101, -108, 90, 93, -47, 67, -125, -90, 23, -88, -32, -87, 46, -102, -10, 83, -77, -66, -105, -62, 126, -10, 125, 54, 0, 84, -60, -78, 52, 14, -21, -17, -97, -66, -104, -68);
    signal scenario_output3 : scenario_type3 :=(-59, -5, 34, -1, 12, -53, 96, 35, -128, -73, 127, 78, -126, -128, 127, -12, 31, 127, -128, 14, 38, 2, -59, 10, 66, -128, 57, 95, -2, 28, -128, -6, 15, -68, 110, -48, 25, 127, -93, -60, 63, 0, 46, 25, -2, 14, -69);
    constant SCENARIO_ADDRESS3 : integer := 49017;    -- This value may arbitrarily change


    constant SCENARIO_LENGTH4 : integer := 24;
    constant SCENARIO_LENGTH_STL4 : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH4, 16));
    type scenario_type4 is array (0 to SCENARIO_LENGTH4-1) of integer;

    signal scenario_config4 : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL4(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL4(7 downto 0))),    -- K2
                                                      0,                                                        -- S
                                                      0, -1, 8, 0, -8, 1, 0, 1, -9, 45, 0, -45, 9, -1           -- C1-C14
                                                      );
    signal scenario_input4 : scenario_type4 := (32, -24, -35,   0, 46, -54, -39, -22, -53, -47,  12, 11,  11, 45, -30, -14, -35, -25, -19, -35, -41, -61, -24, -62);
    signal scenario_output4 : scenario_type4 :=(11,  43, -13, -54, 33,  53, -28,   8,  18, -38, -31,  7, -24, 23,  33,  -1,   7, -11,   5,  10,  15, -12,   3, -10);
 
    constant SCENARIO_ADDRESS4 : integer := 49180;    -- This value may arbitrarily change

    constant SCENARIO_LENGTH5 : integer := 7;
    constant SCENARIO_LENGTH_STL5 : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH5, 16));
    type scenario_type5 is array (0 to SCENARIO_LENGTH5-1) of integer;

    signal scenario_config5 : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL5(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL5(7 downto 0))),    -- K2
                                                      1,                                                        -- S
                                                      0, -1, 8, 0, -8, 1, 0, -128, -128, -128, -128, -128, -128, -128           -- C1-C14
                                                      );
    signal scenario_input5 : scenario_type5 := (127,127,127,127,127,127,127);
    signal scenario_output5 : scenario_type5 :=(-128, -128, -128, -128, -128, -128, -128);
    constant SCENARIO_ADDRESS5 : integer := 49245;  
  
    constant SCENARIO_LENGTH6 : integer := 7;
    constant SCENARIO_LENGTH_STL6 : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH6, 16));
    type scenario_type6 is array (0 to SCENARIO_LENGTH6-1) of integer;

    signal scenario_config6 : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL6(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL6(7 downto 0))),    -- K2
                                                      1,                                                        -- S
                                                      0, -1, 8, 0, -8, 1, 0, -128, -128, -128, -128, -128, -128, -128           -- C1-C14
                                                      );
    signal scenario_input6 : scenario_type6 := (-128, -128, -128, -128, -128, -128, -128);
    signal scenario_output6 : scenario_type6 :=(127,127,127,127,127,127,127);

    constant SCENARIO_ADDRESS6 : integer := 49445;    -- This value may arbitrarily change
  
    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
 
                o_done : out std_logic;
 
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;
 
begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
 
                o_done => tb_done,
 
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );
 
    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;
 
    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
 
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
 
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;
 
        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
 
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;
 
        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';
 
        -- Wait some time for the component to reset...
        wait for 50 ns;
 
        tb_rst <= '0';
        --Start the first run
        memory_control <= '0';  -- Memory controlled by the testbench
 
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock
 
 
        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
 
        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
 
        wait until falling_edge(tb_clk);
 
        memory_control <= '1';  -- Memory controlled by the component
 
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
 
        tb_start <= '1';
 
        --Wait for some time, then reset the component mid elaboration
        for i in 0 to 15 loop
          wait until rising_edge(tb_clk);   
        end loop;
        tb_rst <= '1';
        -- Wait some time for the component to reset...
        wait for 50 ns;
        tb_rst <= '0';
        --Wait for some time, then reset the component mid elaboration (2nd time)
        for i in 0 to 5712 loop
            wait until rising_edge(tb_clk);   
          end loop;
          tb_rst <= '1';
          -- Wait some time for the component to reset...
          wait for 50 ns;
          tb_rst <= '0';
                  
        --Continue with the elaboration
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        wait for 5 ns;
 
        tb_start <= '0';
        
        
        --Start the second run
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS2+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config2(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        for i in 0 to SCENARIO_LENGTH2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS2+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input2(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS2, 16));

        tb_start <= '1';
        
        for i in 0 to 1254 loop
            wait until rising_edge(tb_clk);   
          end loop;
          tb_rst <= '1';
          -- Wait some time for the component to reset...
          wait for 50 ns;
          tb_rst <= '0';
               

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';


        --Start the third run
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS3+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config3(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        for i in 0 to SCENARIO_LENGTH3-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS3+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input3(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS3, 16));

        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

            --RESET
        wait for 50 ns;
 
        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';
 
        -- Wait some time for the component to reset...
        wait for 50 ns;
 
        tb_rst <= '0';


        --Start the forth run
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS4+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config4(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        for i in 0 to SCENARIO_LENGTH4-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS4+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input4(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS4, 16));

        tb_start <= '1';

        for i in 0 to 15 loop
            wait until rising_edge(tb_clk);   
          end loop;
          tb_rst <= '1';
          -- Wait some time for the component to reset...
          wait for 50 ns;
          tb_rst <= '0';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';      

        --start the fifth run
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS5+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config5(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        for i in 0 to SCENARIO_LENGTH5-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS5+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input5(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS5, 16));

        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';            
        
        --start the sixth run
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS6+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config6(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        for i in 0 to SCENARIO_LENGTH6-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS6+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input6(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS6, 16));

        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';            
       
        wait;

    end process;
 
    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin
    
        --Test the first scenario
        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';
 
        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
 
        wait until rising_edge(tb_start);
 
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;
 
        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;
 
        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);
        
        
        --Test the second scenario
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;
 
        for i in 0 to SCENARIO_LENGTH2-1 loop
            assert RAM(SCENARIO_ADDRESS2+17+SCENARIO_LENGTH2+i) = std_logic_vector(to_unsigned(scenario_output2(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH2+i) & " expected= " & integer'image(scenario_output2(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS2+17+SCENARIO_LENGTH2+i)))) severity failure;
        end loop;
 
        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);        

        --Test third scenario
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;
 
        for i in 0 to SCENARIO_LENGTH3-1 loop
            assert RAM(SCENARIO_ADDRESS3+17+SCENARIO_LENGTH3+i) = std_logic_vector(to_unsigned(scenario_output3(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH3+i) & " expected= " & integer'image(scenario_output3(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS3+17+SCENARIO_LENGTH3+i)))) severity failure;
        end loop;
 
        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);        

        --Test forth scenario
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;
 
        for i in 0 to SCENARIO_LENGTH4-1 loop
            assert RAM(SCENARIO_ADDRESS4+17+SCENARIO_LENGTH4+i) = std_logic_vector(to_unsigned(scenario_output4(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH4+i) & " expected= " & integer'image(scenario_output4(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS4+17+SCENARIO_LENGTH4+i)))) severity failure;
        end loop;
 
        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);  

        --Test fifth scenario
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;
 
        for i in 0 to SCENARIO_LENGTH5-1 loop
            assert RAM(SCENARIO_ADDRESS5+17+SCENARIO_LENGTH5+i) = std_logic_vector(to_unsigned(scenario_output5(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH5+i) & " expected= " & integer'image(scenario_output5(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS5+17+SCENARIO_LENGTH5+i)))) severity failure;
        end loop;
 
        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done); 

        --Test sixth scenario
        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;
 
        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;
 
        for i in 0 to SCENARIO_LENGTH6-1 loop
            assert RAM(SCENARIO_ADDRESS6+17+SCENARIO_LENGTH6+i) = std_logic_vector(to_unsigned(scenario_output6(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH6+i) & " expected= " & integer'image(scenario_output6(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS6+17+SCENARIO_LENGTH6+i)))) severity failure;
        end loop;
 
        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);           
  
        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;
 
end architecture;

